module my_chip;
  wire   [15:0] wire_140235384824176;
  wire   [15:0] wire_140235384824176_stb;
  wire   [15:0] wire_140235384824176_ack;
  wire   [15:0] wire_140235384824320;
  wire   [15:0] wire_140235384824320_stb;
  wire   [15:0] wire_140235384824320_ack;
  wire   [15:0] wire_140235384824032;
  wire   [15:0] wire_140235384824032_stb;
  wire   [15:0] wire_140235384824032_ack;
  module 140235384823888_stimulus stimulus(
    wire_140235384824176,
    wire_140235384824176_stb,
    wire_140235384824176_ack);
  module 140235384823960_stimulus stimulus(
    wire_140235384824320,
    wire_140235384824320_stb,
    wire_140235384824320_ack);
  module 140235384716392_adder adder(
    wire_140235384824176,
    wire_140235384824176_stb,
    wire_140235384824176_ack,
    wire_140235384824320,
    wire_140235384824320_stb,
    wire_140235384824320_ack,
    wire_140235384824032,
    wire_140235384824032_stb,
    wire_140235384824032_ack);
  module 140235384717112_response response(
    wire_140235384824032,
    wire_140235384824032_stb,
    wire_140235384824032_ack);
endmodule
