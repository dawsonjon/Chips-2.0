--name: input
--tag: schematic
--output: out1
--source_file: built_in

---Input
---=====
---
---Represents an input to a component in schematix.
