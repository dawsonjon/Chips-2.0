--name: output
--tag: schematic
--input: in_1
--source_file:built_in

---Output
---======
---Used to represent an output from a component in schematix.
