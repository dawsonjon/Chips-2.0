--name: input
--tag: schematic
--output: out1:bits
--source_file: built_in
--parameter: bits:16

---Input
---=====
---
---Represents an input to a component in schematix.
