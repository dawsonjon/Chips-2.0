--name: output
--tag: core
--tag: IO
--input: in_1
--parameter: name : asdfasdfasdf
--source_file:built_in

---Output
---======
---Component Output
