--name: output_16
--tag: schematic
--input: in_1:16
--source_file:built_in

---16-bit Output
---=============
---Used to represent an output from a component in schematix.
