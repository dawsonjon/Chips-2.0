--name: output
--tag: schematic
--input: in_1:bits
--source_file:built_in
--parameter:bits:16

---Output
---======
---Used to represent an output from a component in schematix.
