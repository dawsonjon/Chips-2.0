//name : user_design
//tag : c components
//input : input_checksum:16
//input : input_eth_rx:16
//input : input_rs232_rx:16
//output : output_rs232_tx:16
//output : output_leds:16
//output : output_eth_tx:16
//output : output_checksum:16
//source_file : source/user_design.c
///User_Design
///===========
///
///*Created by C2CHIP*

  
`timescale 1ns/1ps
module user_design(input_checksum,input_eth_rx,input_rs232_rx,input_checksum_stb,input_eth_rx_stb,input_rs232_rx_stb,output_rs232_tx_ack,output_leds_ack,output_eth_tx_ack,output_checksum_ack,clk,rst,output_rs232_tx,output_leds,output_eth_tx,output_checksum,output_rs232_tx_stb,output_leds_stb,output_eth_tx_stb,output_checksum_stb,input_checksum_ack,input_eth_rx_ack,input_rs232_rx_ack);
  input     [15:0] input_checksum;
  input     [15:0] input_eth_rx;
  input     [15:0] input_rs232_rx;
  input     input_checksum_stb;
  input     input_eth_rx_stb;
  input     input_rs232_rx_stb;
  input     output_rs232_tx_ack;
  input     output_leds_ack;
  input     output_eth_tx_ack;
  input     output_checksum_ack;
  input     clk;
  input     rst;
  output    [15:0] output_rs232_tx;
  output    [15:0] output_leds;
  output    [15:0] output_eth_tx;
  output    [15:0] output_checksum;
  output    output_rs232_tx_stb;
  output    output_leds_stb;
  output    output_eth_tx_stb;
  output    output_checksum_stb;
  output    input_checksum_ack;
  output    input_eth_rx_ack;
  output    input_rs232_rx_ack;
  reg       [15:0] timer;
  reg       [9:0] program_counter;
  reg       [15:0] address;
  reg       [15:0] data_out;
  reg       [15:0] data_in;
  reg       write_enable;
  reg       [15:0] register_0;
  reg       [15:0] register_1;
  reg       [15:0] register_2;
  reg       [15:0] register_3;
  reg       [15:0] register_4;
  reg       [15:0] register_5;
  reg       [15:0] register_6;
  reg       [15:0] register_7;
  reg       [15:0] register_8;
  reg       [15:0] register_9;
  reg       [15:0] register_10;
  reg       [15:0] register_11;
  reg       [15:0] register_12;
  reg       [15:0] register_13;
  reg       [15:0] register_14;
  reg       [15:0] register_15;
  reg       [15:0] register_16;
  reg       [15:0] register_17;
  reg       [15:0] register_18;
  reg       [15:0] register_19;
  reg       [15:0] register_20;
  reg       [15:0] register_21;
  reg       [15:0] register_22;
  reg       [15:0] register_23;
  reg       [15:0] register_24;
  reg       [15:0] register_25;
  reg       [15:0] register_26;
  reg       [15:0] register_27;
  reg       [15:0] register_28;
  reg       [15:0] register_29;
  reg       [15:0] register_30;
  reg       [15:0] register_31;
  reg       [15:0] register_32;
  reg       [15:0] register_33;
  reg       [15:0] register_34;
  reg       [15:0] register_35;
  reg       [15:0] register_36;
  reg       [15:0] register_37;
  reg       [15:0] register_38;
  reg       [15:0] register_39;
  reg       [15:0] register_40;
  reg       [15:0] register_41;
  reg       [15:0] register_42;
  reg       [15:0] register_43;
  reg       [15:0] register_44;
  reg       [15:0] register_45;
  reg       [15:0] register_46;
  reg       [15:0] register_47;
  reg       [15:0] register_48;
  reg       [15:0] register_49;
  reg       [15:0] register_50;
  reg       [15:0] register_51;
  reg       [15:0] register_52;
  reg       [15:0] register_53;
  reg       [15:0] register_54;
  reg       [15:0] register_55;
  reg       [15:0] register_56;
  reg       [15:0] register_57;
  reg       [15:0] register_58;
  reg       [15:0] register_59;
  reg       [15:0] register_60;
  reg       [15:0] register_61;
  reg       [15:0] register_62;
  reg       [15:0] register_63;
  reg       [15:0] register_64;
  reg       [15:0] register_65;
  reg       [15:0] register_66;
  reg       [15:0] register_67;
  reg       [15:0] register_68;
  reg       [15:0] register_69;
  reg       [15:0] register_70;
  reg       [15:0] register_71;
  reg       [15:0] register_72;
  reg       [15:0] register_73;
  reg       [15:0] register_74;
  reg       [15:0] register_75;
  reg       [15:0] register_76;
  reg       [15:0] register_77;
  reg       [15:0] register_78;
  reg       [15:0] register_79;
  reg       [15:0] register_80;
  reg       [15:0] register_81;
  reg       [15:0] register_82;
  reg       [15:0] register_83;
  reg       [15:0] register_84;
  reg       [15:0] register_85;
  reg       [15:0] register_86;
  reg       [15:0] register_87;
  reg       [15:0] register_88;
  reg       [15:0] register_89;
  reg       [15:0] register_90;
  reg       [15:0] register_91;
  reg       [15:0] register_92;
  reg       [15:0] register_93;
  reg       [15:0] register_94;
  reg       [15:0] register_95;
  reg       [15:0] register_96;
  reg       [15:0] register_97;
  reg       [15:0] register_98;
  reg       [15:0] register_99;
  reg       [15:0] register_100;
  reg       [15:0] register_101;
  reg       [15:0] register_102;
  reg       [15:0] register_103;
  reg       [15:0] register_104;
  reg       [15:0] register_105;
  reg       [15:0] register_106;
  reg       [15:0] register_107;
  reg       [15:0] register_108;
  reg       [15:0] register_109;
  reg       [15:0] register_110;
  reg       [15:0] register_111;
  reg       [15:0] register_112;
  reg       [15:0] register_113;
  reg       [15:0] register_114;
  reg       [15:0] register_115;
  reg       [15:0] register_116;
  reg       [15:0] register_117;
  reg       [15:0] register_118;
  reg       [15:0] register_119;
  reg       [15:0] register_120;
  reg       [15:0] register_121;
  reg       [15:0] register_122;
  reg       [15:0] register_123;
  reg       [15:0] register_124;
  reg       [15:0] register_125;
  reg       [15:0] register_126;
  reg       [15:0] register_127;
  reg       [15:0] register_128;
  reg       [15:0] register_129;
  reg       [15:0] register_130;
  reg       [15:0] register_131;
  reg       [15:0] register_132;
  reg       [15:0] register_133;
  reg       [15:0] register_134;
  reg       [15:0] register_135;
  reg       [15:0] register_136;
  reg       [15:0] register_137;
  reg       [15:0] register_138;
  reg       [15:0] register_139;
  reg       [15:0] register_140;
  reg       [15:0] register_141;
  reg       [15:0] register_142;
  reg       [15:0] register_143;
  reg       [15:0] register_144;
  reg       [15:0] register_145;
  reg       [15:0] register_146;
  reg       [15:0] register_147;
  reg       [15:0] register_148;
  reg       [15:0] register_149;
  reg       [15:0] register_150;
  reg       [15:0] register_151;
  reg       [15:0] register_152;
  reg       [15:0] register_153;
  reg       [15:0] register_154;
  reg       [15:0] register_155;
  reg       [15:0] register_156;
  reg       [15:0] register_157;
  reg       [15:0] register_158;
  reg       [15:0] register_159;
  reg       [15:0] register_160;
  reg       [15:0] register_161;
  reg       [15:0] register_162;
  reg       [15:0] register_163;
  reg       [15:0] register_164;
  reg       [15:0] register_165;
  reg       [15:0] register_166;
  reg       [15:0] register_167;
  reg       [15:0] register_168;
  reg       [15:0] register_169;
  reg       [15:0] register_170;
  reg       [15:0] register_171;
  reg       [15:0] register_172;
  reg       [15:0] register_173;
  reg       [15:0] s_output_rs232_tx_stb;
  reg       [15:0] s_output_leds_stb;
  reg       [15:0] s_output_eth_tx_stb;
  reg       [15:0] s_output_checksum_stb;
  reg       [15:0] s_output_rs232_tx;
  reg       [15:0] s_output_leds;
  reg       [15:0] s_output_eth_tx;
  reg       [15:0] s_output_checksum;
  reg       [15:0] s_input_checksum_ack;
  reg       [15:0] s_input_eth_rx_ack;
  reg       [15:0] s_input_rs232_rx_ack;
  reg [15:0] memory [3088:0];

  //////////////////////////////////////////////////////////////////////////////
  // MEMORY INITIALIZATION                                                      
  //                                                                            
  // In order to reduce program size, array contents have been stored into      
  // memory at initialization. In an FPGA, this will result in the memory being 
  // initialized when the FPGA configures.                                      
  // Memory will not be re-initialized at reset.                                
  // Dissable this behaviour using the no_initialize_memory switch              
  
  initial
  begin
    memory[16'd512] = 16'd112;
    memory[16'd513] = 16'd117;
    memory[16'd514] = 16'd116;
    memory[16'd515] = 16'd95;
    memory[16'd516] = 16'd101;
    memory[16'd517] = 16'd116;
    memory[16'd518] = 16'd104;
    memory[16'd519] = 16'd10;
    memory[16'd520] = 16'd0;
    memory[16'd521] = 16'd103;
    memory[16'd522] = 16'd101;
    memory[16'd523] = 16'd116;
    memory[16'd524] = 16'd95;
    memory[16'd525] = 16'd101;
    memory[16'd526] = 16'd116;
    memory[16'd527] = 16'd104;
    memory[16'd528] = 16'd10;
    memory[16'd529] = 16'd0;
    memory[16'd530] = 16'd114;
    memory[16'd531] = 16'd101;
    memory[16'd532] = 16'd97;
    memory[16'd533] = 16'd100;
    memory[16'd534] = 16'd105;
    memory[16'd535] = 16'd110;
    memory[16'd536] = 16'd103;
    memory[16'd537] = 16'd32;
    memory[16'd538] = 16'd98;
    memory[16'd539] = 16'd121;
    memory[16'd540] = 16'd116;
    memory[16'd541] = 16'd101;
    memory[16'd542] = 16'd115;
    memory[16'd543] = 16'd58;
    memory[16'd544] = 16'd32;
    memory[16'd545] = 16'd0;
    memory[16'd546] = 16'd10;
    memory[16'd547] = 16'd0;
    memory[16'd548] = 16'd100;
    memory[16'd549] = 16'd111;
    memory[16'd550] = 16'd110;
    memory[16'd551] = 16'd101;
    memory[16'd552] = 16'd10;
    memory[16'd553] = 16'd0;
    memory[16'd554] = 16'd10;
    memory[16'd555] = 16'd0;
    memory[16'd556] = 16'd10;
    memory[16'd557] = 16'd0;
    memory[16'd558] = 16'd10;
    memory[16'd559] = 16'd0;
    memory[16'd560] = 16'd109;
    memory[16'd561] = 16'd97;
    memory[16'd562] = 16'd99;
    memory[16'd563] = 16'd32;
    memory[16'd564] = 16'd103;
    memory[16'd565] = 16'd111;
    memory[16'd566] = 16'd111;
    memory[16'd567] = 16'd100;
    memory[16'd568] = 16'd10;
    memory[16'd569] = 16'd0;
    memory[16'd570] = 16'd97;
    memory[16'd571] = 16'd114;
    memory[16'd572] = 16'd112;
    memory[16'd573] = 16'd10;
    memory[16'd574] = 16'd0;
    memory[16'd671] = 16'd99;
    memory[16'd672] = 16'd97;
    memory[16'd673] = 16'd99;
    memory[16'd674] = 16'd104;
    memory[16'd675] = 16'd101;
    memory[16'd676] = 16'd32;
    memory[16'd677] = 16'd104;
    memory[16'd678] = 16'd105;
    memory[16'd679] = 16'd116;
    memory[16'd680] = 16'd10;
    memory[16'd681] = 16'd0;
    memory[16'd682] = 16'd99;
    memory[16'd683] = 16'd97;
    memory[16'd684] = 16'd99;
    memory[16'd685] = 16'd104;
    memory[16'd686] = 16'd101;
    memory[16'd687] = 16'd32;
    memory[16'd688] = 16'd109;
    memory[16'd689] = 16'd105;
    memory[16'd690] = 16'd115;
    memory[16'd691] = 16'd115;
    memory[16'd692] = 16'd10;
    memory[16'd693] = 16'd0;
    memory[16'd694] = 16'd97;
    memory[16'd695] = 16'd114;
    memory[16'd696] = 16'd112;
    memory[16'd697] = 16'd32;
    memory[16'd698] = 16'd114;
    memory[16'd699] = 16'd101;
    memory[16'd700] = 16'd113;
    memory[16'd701] = 16'd117;
    memory[16'd702] = 16'd101;
    memory[16'd703] = 16'd115;
    memory[16'd704] = 16'd116;
    memory[16'd705] = 16'd10;
    memory[16'd706] = 16'd0;
    memory[16'd707] = 16'd103;
    memory[16'd708] = 16'd111;
    memory[16'd709] = 16'd116;
    memory[16'd710] = 16'd95;
    memory[16'd711] = 16'd112;
    memory[16'd712] = 16'd97;
    memory[16'd713] = 16'd99;
    memory[16'd714] = 16'd107;
    memory[16'd715] = 16'd101;
    memory[16'd716] = 16'd116;
    memory[16'd717] = 16'd10;
    memory[16'd718] = 16'd0;
    memory[16'd719] = 16'd97;
    memory[16'd720] = 16'd114;
    memory[16'd721] = 16'd112;
    memory[16'd722] = 16'd32;
    memory[16'd723] = 16'd114;
    memory[16'd724] = 16'd101;
    memory[16'd725] = 16'd115;
    memory[16'd726] = 16'd112;
    memory[16'd727] = 16'd111;
    memory[16'd728] = 16'd110;
    memory[16'd729] = 16'd115;
    memory[16'd730] = 16'd101;
    memory[16'd731] = 16'd10;
    memory[16'd732] = 16'd0;
    memory[16'd733] = 16'd117;
    memory[16'd734] = 16'd112;
    memory[16'd735] = 16'd100;
    memory[16'd736] = 16'd97;
    memory[16'd737] = 16'd116;
    memory[16'd738] = 16'd105;
    memory[16'd739] = 16'd110;
    memory[16'd740] = 16'd103;
    memory[16'd741] = 16'd32;
    memory[16'd742] = 16'd99;
    memory[16'd743] = 16'd97;
    memory[16'd744] = 16'd99;
    memory[16'd745] = 16'd104;
    memory[16'd746] = 16'd101;
    memory[16'd747] = 16'd10;
    memory[16'd748] = 16'd0;
    memory[16'd749] = 16'd112;
    memory[16'd750] = 16'd117;
    memory[16'd751] = 16'd116;
    memory[16'd752] = 16'd95;
    memory[16'd753] = 16'd105;
    memory[16'd754] = 16'd112;
    memory[16'd755] = 16'd10;
    memory[16'd756] = 16'd0;
    memory[16'd757] = 16'd103;
    memory[16'd758] = 16'd101;
    memory[16'd759] = 16'd116;
    memory[16'd760] = 16'd95;
    memory[16'd761] = 16'd105;
    memory[16'd762] = 16'd112;
    memory[16'd763] = 16'd10;
    memory[16'd764] = 16'd0;
    memory[16'd765] = 16'd105;
    memory[16'd766] = 16'd112;
    memory[16'd767] = 16'd10;
    memory[16'd768] = 16'd0;
    memory[16'd769] = 16'd105;
    memory[16'd770] = 16'd112;
    memory[16'd771] = 16'd32;
    memory[16'd772] = 16'd97;
    memory[16'd773] = 16'd100;
    memory[16'd774] = 16'd100;
    memory[16'd775] = 16'd114;
    memory[16'd776] = 16'd101;
    memory[16'd777] = 16'd115;
    memory[16'd778] = 16'd115;
    memory[16'd779] = 16'd32;
    memory[16'd780] = 16'd103;
    memory[16'd781] = 16'd111;
    memory[16'd782] = 16'd111;
    memory[16'd783] = 16'd100;
    memory[16'd784] = 16'd10;
    memory[16'd785] = 16'd0;
    memory[16'd786] = 16'd105;
    memory[16'd787] = 16'd99;
    memory[16'd788] = 16'd109;
    memory[16'd789] = 16'd112;
    memory[16'd790] = 16'd10;
    memory[16'd791] = 16'd0;
    memory[16'd792] = 16'd112;
    memory[16'd793] = 16'd105;
    memory[16'd794] = 16'd110;
    memory[16'd795] = 16'd103;
    memory[16'd796] = 16'd95;
    memory[16'd797] = 16'd114;
    memory[16'd798] = 16'd101;
    memory[16'd799] = 16'd113;
    memory[16'd800] = 16'd117;
    memory[16'd801] = 16'd101;
    memory[16'd802] = 16'd115;
    memory[16'd803] = 16'd116;
    memory[16'd804] = 16'd10;
    memory[16'd805] = 16'd0;
    memory[16'd806] = 16'd111;
    memory[16'd807] = 16'd116;
    memory[16'd808] = 16'd104;
    memory[16'd809] = 16'd101;
    memory[16'd810] = 16'd114;
    memory[16'd811] = 16'd0;
    memory[16'd812] = 16'd112;
    memory[16'd813] = 16'd117;
    memory[16'd814] = 16'd116;
    memory[16'd815] = 16'd32;
    memory[16'd816] = 16'd116;
    memory[16'd817] = 16'd99;
    memory[16'd818] = 16'd112;
    memory[16'd819] = 16'd10;
    memory[16'd820] = 16'd0;
    memory[16'd821] = 16'd103;
    memory[16'd822] = 16'd101;
    memory[16'd823] = 16'd116;
    memory[16'd824] = 16'd32;
    memory[16'd825] = 16'd116;
    memory[16'd826] = 16'd99;
    memory[16'd827] = 16'd112;
    memory[16'd828] = 16'd10;
    memory[16'd829] = 16'd0;
    memory[16'd830] = 16'd115;
    memory[16'd831] = 16'd111;
    memory[16'd832] = 16'd117;
    memory[16'd833] = 16'd114;
    memory[16'd834] = 16'd99;
    memory[16'd835] = 16'd101;
    memory[16'd836] = 16'd58;
    memory[16'd837] = 16'd32;
    memory[16'd838] = 16'd0;
    memory[16'd839] = 16'd10;
    memory[16'd840] = 16'd0;
    memory[16'd841] = 16'd100;
    memory[16'd842] = 16'd101;
    memory[16'd843] = 16'd115;
    memory[16'd844] = 16'd116;
    memory[16'd845] = 16'd58;
    memory[16'd846] = 16'd32;
    memory[16'd847] = 16'd0;
    memory[16'd848] = 16'd10;
    memory[16'd849] = 16'd0;
    memory[16'd850] = 16'd115;
    memory[16'd851] = 16'd101;
    memory[16'd852] = 16'd113;
    memory[16'd853] = 16'd95;
    memory[16'd854] = 16'd104;
    memory[16'd855] = 16'd105;
    memory[16'd856] = 16'd58;
    memory[16'd857] = 16'd32;
    memory[16'd858] = 16'd0;
    memory[16'd859] = 16'd10;
    memory[16'd860] = 16'd0;
    memory[16'd861] = 16'd115;
    memory[16'd862] = 16'd101;
    memory[16'd863] = 16'd113;
    memory[16'd864] = 16'd95;
    memory[16'd865] = 16'd108;
    memory[16'd866] = 16'd111;
    memory[16'd867] = 16'd58;
    memory[16'd868] = 16'd32;
    memory[16'd869] = 16'd0;
    memory[16'd870] = 16'd10;
    memory[16'd871] = 16'd0;
    memory[16'd872] = 16'd97;
    memory[16'd873] = 16'd99;
    memory[16'd874] = 16'd107;
    memory[16'd875] = 16'd95;
    memory[16'd876] = 16'd104;
    memory[16'd877] = 16'd105;
    memory[16'd878] = 16'd58;
    memory[16'd879] = 16'd32;
    memory[16'd880] = 16'd0;
    memory[16'd881] = 16'd10;
    memory[16'd882] = 16'd0;
    memory[16'd883] = 16'd97;
    memory[16'd884] = 16'd99;
    memory[16'd885] = 16'd107;
    memory[16'd886] = 16'd95;
    memory[16'd887] = 16'd108;
    memory[16'd888] = 16'd111;
    memory[16'd889] = 16'd58;
    memory[16'd890] = 16'd32;
    memory[16'd891] = 16'd0;
    memory[16'd892] = 16'd10;
    memory[16'd893] = 16'd0;
    memory[16'd894] = 16'd119;
    memory[16'd895] = 16'd105;
    memory[16'd896] = 16'd110;
    memory[16'd897] = 16'd100;
    memory[16'd898] = 16'd111;
    memory[16'd899] = 16'd119;
    memory[16'd900] = 16'd58;
    memory[16'd901] = 16'd32;
    memory[16'd902] = 16'd0;
    memory[16'd903] = 16'd10;
    memory[16'd904] = 16'd0;
    memory[16'd905] = 16'd102;
    memory[16'd906] = 16'd108;
    memory[16'd907] = 16'd97;
    memory[16'd908] = 16'd103;
    memory[16'd909] = 16'd115;
    memory[16'd910] = 16'd58;
    memory[16'd911] = 16'd32;
    memory[16'd912] = 16'd0;
    memory[16'd913] = 16'd10;
    memory[16'd914] = 16'd0;
    memory[16'd2963] = 16'd10;
    memory[16'd2964] = 16'd69;
    memory[16'd2965] = 16'd116;
    memory[16'd2966] = 16'd104;
    memory[16'd2967] = 16'd101;
    memory[16'd2968] = 16'd114;
    memory[16'd2969] = 16'd110;
    memory[16'd2970] = 16'd101;
    memory[16'd2971] = 16'd116;
    memory[16'd2972] = 16'd32;
    memory[16'd2973] = 16'd77;
    memory[16'd2974] = 16'd111;
    memory[16'd2975] = 16'd110;
    memory[16'd2976] = 16'd105;
    memory[16'd2977] = 16'd116;
    memory[16'd2978] = 16'd111;
    memory[16'd2979] = 16'd114;
    memory[16'd2980] = 16'd10;
    memory[16'd2981] = 16'd0;
    memory[16'd2982] = 16'd119;
    memory[16'd2983] = 16'd97;
    memory[16'd2984] = 16'd105;
    memory[16'd2985] = 16'd116;
    memory[16'd2986] = 16'd105;
    memory[16'd2987] = 16'd110;
    memory[16'd2988] = 16'd103;
    memory[16'd2989] = 16'd32;
    memory[16'd2990] = 16'd102;
    memory[16'd2991] = 16'd111;
    memory[16'd2992] = 16'd114;
    memory[16'd2993] = 16'd32;
    memory[16'd2994] = 16'd99;
    memory[16'd2995] = 16'd111;
    memory[16'd2996] = 16'd110;
    memory[16'd2997] = 16'd110;
    memory[16'd2998] = 16'd101;
    memory[16'd2999] = 16'd99;
    memory[16'd3000] = 16'd116;
    memory[16'd3001] = 16'd105;
    memory[16'd3002] = 16'd111;
    memory[16'd3003] = 16'd110;
    memory[16'd3004] = 16'd10;
    memory[16'd3005] = 16'd0;
    memory[16'd3006] = 16'd105;
    memory[16'd3007] = 16'd110;
    memory[16'd3008] = 16'd99;
    memory[16'd3009] = 16'd111;
    memory[16'd3010] = 16'd109;
    memory[16'd3011] = 16'd109;
    memory[16'd3012] = 16'd105;
    memory[16'd3013] = 16'd110;
    memory[16'd3014] = 16'd103;
    memory[16'd3015] = 16'd32;
    memory[16'd3016] = 16'd99;
    memory[16'd3017] = 16'd111;
    memory[16'd3018] = 16'd110;
    memory[16'd3019] = 16'd110;
    memory[16'd3020] = 16'd101;
    memory[16'd3021] = 16'd99;
    memory[16'd3022] = 16'd116;
    memory[16'd3023] = 16'd105;
    memory[16'd3024] = 16'd111;
    memory[16'd3025] = 16'd110;
    memory[16'd3026] = 16'd32;
    memory[16'd3027] = 16'd102;
    memory[16'd3028] = 16'd114;
    memory[16'd3029] = 16'd111;
    memory[16'd3030] = 16'd109;
    memory[16'd3031] = 16'd58;
    memory[16'd3032] = 16'd32;
    memory[16'd3033] = 16'd0;
    memory[16'd3034] = 16'd10;
    memory[16'd3035] = 16'd0;
    memory[16'd3036] = 16'd119;
    memory[16'd3037] = 16'd97;
    memory[16'd3038] = 16'd105;
    memory[16'd3039] = 16'd116;
    memory[16'd3040] = 16'd105;
    memory[16'd3041] = 16'd110;
    memory[16'd3042] = 16'd103;
    memory[16'd3043] = 16'd32;
    memory[16'd3044] = 16'd102;
    memory[16'd3045] = 16'd111;
    memory[16'd3046] = 16'd114;
    memory[16'd3047] = 16'd32;
    memory[16'd3048] = 16'd97;
    memory[16'd3049] = 16'd99;
    memory[16'd3050] = 16'd107;
    memory[16'd3051] = 16'd110;
    memory[16'd3052] = 16'd111;
    memory[16'd3053] = 16'd119;
    memory[16'd3054] = 16'd108;
    memory[16'd3055] = 16'd101;
    memory[16'd3056] = 16'd100;
    memory[16'd3057] = 16'd103;
    memory[16'd3058] = 16'd101;
    memory[16'd3059] = 16'd109;
    memory[16'd3060] = 16'd101;
    memory[16'd3061] = 16'd110;
    memory[16'd3062] = 16'd116;
    memory[16'd3063] = 16'd10;
    memory[16'd3064] = 16'd0;
    memory[16'd3065] = 16'd99;
    memory[16'd3066] = 16'd111;
    memory[16'd3067] = 16'd110;
    memory[16'd3068] = 16'd110;
    memory[16'd3069] = 16'd101;
    memory[16'd3070] = 16'd99;
    memory[16'd3071] = 16'd116;
    memory[16'd3072] = 16'd105;
    memory[16'd3073] = 16'd111;
    memory[16'd3074] = 16'd110;
    memory[16'd3075] = 16'd32;
    memory[16'd3076] = 16'd101;
    memory[16'd3077] = 16'd115;
    memory[16'd3078] = 16'd116;
    memory[16'd3079] = 16'd97;
    memory[16'd3080] = 16'd98;
    memory[16'd3081] = 16'd108;
    memory[16'd3082] = 16'd105;
    memory[16'd3083] = 16'd115;
    memory[16'd3084] = 16'd104;
    memory[16'd3085] = 16'd101;
    memory[16'd3086] = 16'd100;
    memory[16'd3087] = 16'd10;
    memory[16'd3088] = 16'd0;
  end


  //////////////////////////////////////////////////////////////////////////////
  // FSM IMPLEMENTAION OF C PROCESS                                             
  //                                                                            
  // This section of the file contains a Finite State Machine (FSM) implementing
  // the C process. In general execution is sequential, but the compiler will   
  // attempt to execute instructions in parallel if the instruction dependencies
  // allow. Further concurrency can be achieved by executing multiple C         
  // processes concurrently within the device.                                  
  
  always @(posedge clk)
  begin

    if (write_enable == 1'b1) begin
      memory[address] <= data_in;
    end

    data_out <= memory[address];
    write_enable <= 1'b0;
    program_counter <= program_counter + 1;
    timer <= 16'h0000;

    case(program_counter)

      16'd0:
      begin
        register_0 <= 16'd1;
        register_1 <= 16'd515;
        register_2 <= 16'd1029;
        register_3 <= 16'd49320;
        register_4 <= 16'd257;
        register_5 <= 16'd23;
        register_6 <= 16'd0;
        register_43 <= 16'd575;
        register_44 <= 16'd591;
        register_45 <= 16'd607;
        register_46 <= 16'd623;
        register_47 <= 16'd639;
        register_48 <= 16'd0;
        register_92 <= 16'd0;
        register_93 <= 16'd0;
        register_94 <= 16'd0;
        register_95 <= 16'd0;
        register_96 <= 16'd0;
        register_97 <= 16'd0;
        register_98 <= 16'd0;
        register_99 <= 16'd0;
        register_100 <= 16'd255;
        register_101 <= 16'd0;
        register_102 <= 16'd0;
        register_103 <= 16'd0;
        register_104 <= 16'd0;
        register_105 <= 16'd0;
        register_106 <= 16'd0;
        register_107 <= 16'd0;
        register_108 <= 16'd0;
        register_109 <= 16'd0;
        register_110 <= 16'd0;
        register_111 <= 16'd0;
        register_112 <= 16'd0;
        register_113 <= 16'd0;
        register_114 <= 16'd0;
        register_115 <= 16'd0;
        register_116 <= 16'd0;
        register_117 <= 16'd0;
        register_118 <= 16'd0;
        register_119 <= 16'd0;
        program_counter <= 16'd924;
        register_157 <= 16'd1;
      end

      16'd1:
      begin
        program_counter <= program_counter;
      end

      16'd2:
      begin
        register_10 <= 16'd0;
      end

      16'd3:
      begin
        register_172 <= register_10;
      end

      16'd4:
      begin
        register_172 <= $signed(register_172) + $signed(register_9);
      end

      16'd5:
      begin
        address <= register_172;
      end

      16'd6:
      begin
        register_172 <= data_out;
      end

      16'd7:
      begin
        register_172 <= data_out;
      end

      16'd8:
      begin
        register_172 <= $signed(register_172) != $signed(16'd0);
      end

      16'd9:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 19;
      end

      16'd10:
      begin
        register_172 <= register_10;
      end

      16'd11:
      begin
        register_172 <= $signed(register_172) + $signed(register_9);
      end

      16'd12:
      begin
        address <= register_172;
      end

      16'd13:
      begin
        register_172 <= data_out;
      end

      16'd14:
      begin
        register_172 <= data_out;
      end

      16'd15:
      begin
        s_output_rs232_tx <= register_172;
        program_counter <= 15;
        s_output_rs232_tx_stb <= 1'b1;
        if (s_output_rs232_tx_stb == 1'b1 && output_rs232_tx_ack == 1'b1) begin
          s_output_rs232_tx_stb <= 1'b0;
          program_counter <= 16;
        end
      end

      16'd16:
      begin
        register_172 <= register_10;
      end

      16'd17:
      begin
        register_172 <= $signed(register_172) + $signed(16'd1);
      end

      16'd18:
      begin
        register_10 <= register_172;
        program_counter <= 16'd20;
      end

      16'd19:
      begin
        program_counter <= 16'd21;
      end

      16'd20:
      begin
        program_counter <= 16'd3;
      end

      16'd21:
      begin
        register_8 <= 16'd0;
        program_counter <= register_7;
      end

      16'd22:
      begin
        register_172 <= register_13;
      end

      16'd23:
      begin
        register_172 <= $signed(register_172) > $signed(16'd9);
      end

      16'd24:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 28;
      end

      16'd25:
      begin
        register_12 <= register_13;
      end

      16'd26:
      begin
        register_12 <= $signed(register_12) + $signed(16'd87);
        program_counter <= register_11;
      end

      16'd27:
      begin
        program_counter <= 16'd28;
      end

      16'd28:
      begin
        register_12 <= register_13;
      end

      16'd29:
      begin
        register_12 <= $signed(register_12) + $signed(16'd48);
        program_counter <= register_11;
      end

      16'd30:
      begin
        register_13 <= register_16;
      end

      16'd31:
      begin
        register_13 <= $signed(register_13) >>> $signed(16'd12);
      end

      16'd32:
      begin
        register_13 <= $signed(register_13) & $signed(16'd15);
        program_counter <= 16'd22;
        register_11 <= 16'd33;
      end

      16'd33:
      begin
        register_172 <= register_12;
      end

      16'd34:
      begin
        s_output_rs232_tx <= register_172;
        program_counter <= 34;
        s_output_rs232_tx_stb <= 1'b1;
        if (s_output_rs232_tx_stb == 1'b1 && output_rs232_tx_ack == 1'b1) begin
          s_output_rs232_tx_stb <= 1'b0;
          program_counter <= 35;
        end
      end

      16'd35:
      begin
        register_13 <= register_16;
      end

      16'd36:
      begin
        register_13 <= $signed(register_13) >>> $signed(16'd8);
      end

      16'd37:
      begin
        register_13 <= $signed(register_13) & $signed(16'd15);
        program_counter <= 16'd22;
        register_11 <= 16'd38;
      end

      16'd38:
      begin
        register_172 <= register_12;
      end

      16'd39:
      begin
        s_output_rs232_tx <= register_172;
        program_counter <= 39;
        s_output_rs232_tx_stb <= 1'b1;
        if (s_output_rs232_tx_stb == 1'b1 && output_rs232_tx_ack == 1'b1) begin
          s_output_rs232_tx_stb <= 1'b0;
          program_counter <= 40;
        end
      end

      16'd40:
      begin
        register_172 <= 16'd32;
      end

      16'd41:
      begin
        s_output_rs232_tx <= register_172;
        program_counter <= 41;
        s_output_rs232_tx_stb <= 1'b1;
        if (s_output_rs232_tx_stb == 1'b1 && output_rs232_tx_ack == 1'b1) begin
          s_output_rs232_tx_stb <= 1'b0;
          program_counter <= 42;
        end
      end

      16'd42:
      begin
        register_13 <= register_16;
      end

      16'd43:
      begin
        register_13 <= $signed(register_13) >>> $signed(16'd4);
      end

      16'd44:
      begin
        register_13 <= $signed(register_13) & $signed(16'd15);
        program_counter <= 16'd22;
        register_11 <= 16'd45;
      end

      16'd45:
      begin
        register_172 <= register_12;
      end

      16'd46:
      begin
        s_output_rs232_tx <= register_172;
        program_counter <= 46;
        s_output_rs232_tx_stb <= 1'b1;
        if (s_output_rs232_tx_stb == 1'b1 && output_rs232_tx_ack == 1'b1) begin
          s_output_rs232_tx_stb <= 1'b0;
          program_counter <= 47;
        end
      end

      16'd47:
      begin
        register_13 <= register_16;
      end

      16'd48:
      begin
        register_13 <= $signed(register_13) & $signed(16'd15);
        program_counter <= 16'd22;
        register_11 <= 16'd49;
      end

      16'd49:
      begin
        register_172 <= register_12;
      end

      16'd50:
      begin
        s_output_rs232_tx <= register_172;
        program_counter <= 50;
        s_output_rs232_tx_stb <= 1'b1;
        if (s_output_rs232_tx_stb == 1'b1 && output_rs232_tx_ack == 1'b1) begin
          s_output_rs232_tx_stb <= 1'b0;
          program_counter <= 51;
        end
      end

      16'd51:
      begin
        register_172 <= 16'd32;
      end

      16'd52:
      begin
        s_output_rs232_tx <= register_172;
        program_counter <= 52;
        s_output_rs232_tx_stb <= 1'b1;
        if (s_output_rs232_tx_stb == 1'b1 && output_rs232_tx_ack == 1'b1) begin
          s_output_rs232_tx_stb <= 1'b0;
          program_counter <= 53;
        end
      end

      16'd53:
      begin
        register_15 <= 16'd0;
        program_counter <= register_14;
      end

      16'd54:
      begin
        register_25 <= 16'd0;
        register_26 <= 16'd0;
        register_27 <= 16'd512;
      end

      16'd55:
      begin
        register_9 <= register_27;
        program_counter <= 16'd2;
        register_7 <= 16'd56;
      end

      16'd56:
      begin
        register_172 <= register_8;
        register_173 <= 16'd0;
      end

      16'd57:
      begin
        register_172 <= register_21;
        register_173 <= $signed(register_173) + $signed(register_19);
      end

      16'd58:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_22;
        register_173 <= 16'd1;
      end

      16'd59:
      begin
        register_173 <= $signed(register_173) + $signed(register_19);
      end

      16'd60:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_23;
        register_173 <= 16'd2;
      end

      16'd61:
      begin
        register_173 <= $signed(register_173) + $signed(register_19);
      end

      16'd62:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_0;
        register_173 <= 16'd3;
      end

      16'd63:
      begin
        register_173 <= $signed(register_173) + $signed(register_19);
      end

      16'd64:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_1;
        register_173 <= 16'd4;
      end

      16'd65:
      begin
        register_173 <= $signed(register_173) + $signed(register_19);
      end

      16'd66:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_2;
        register_173 <= 16'd5;
      end

      16'd67:
      begin
        register_173 <= $signed(register_173) + $signed(register_19);
      end

      16'd68:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_24;
        register_173 <= 16'd6;
      end

      16'd69:
      begin
        register_173 <= $signed(register_173) + $signed(register_19);
      end

      16'd70:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_20;
      end

      16'd71:
      begin
        s_output_eth_tx <= register_172;
        program_counter <= 71;
        s_output_eth_tx_stb <= 1'b1;
        if (s_output_eth_tx_stb == 1'b1 && output_eth_tx_ack == 1'b1) begin
          s_output_eth_tx_stb <= 1'b0;
          program_counter <= 72;
        end
      end

      16'd72:
      begin
        register_172 <= 16'd0;
      end

      16'd73:
      begin
        register_26 <= register_172;
        register_172 <= 16'd0;
      end

      16'd74:
      begin
        register_25 <= register_172;
      end

      16'd75:
      begin
        register_172 <= register_25;
        register_173 <= register_20;
      end

      16'd76:
      begin
        register_172 <= $signed(register_172) < $signed(register_173);
      end

      16'd77:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 90;
      end

      16'd78:
      begin
        register_172 <= register_26;
      end

      16'd79:
      begin
        register_172 <= $signed(register_172) + $signed(register_19);
      end

      16'd80:
      begin
        address <= register_172;
      end

      16'd81:
      begin
        register_172 <= data_out;
      end

      16'd82:
      begin
        register_172 <= data_out;
      end

      16'd83:
      begin
        s_output_eth_tx <= register_172;
        program_counter <= 83;
        s_output_eth_tx_stb <= 1'b1;
        if (s_output_eth_tx_stb == 1'b1 && output_eth_tx_ack == 1'b1) begin
          s_output_eth_tx_stb <= 1'b0;
          program_counter <= 84;
        end
      end

      16'd84:
      begin
        register_172 <= register_26;
      end

      16'd85:
      begin
        register_172 <= $signed(register_172) + $signed(16'd1);
      end

      16'd86:
      begin
        register_26 <= register_172;
      end

      16'd87:
      begin
        register_172 <= register_25;
      end

      16'd88:
      begin
        register_172 <= $signed(register_172) + $signed(16'd2);
      end

      16'd89:
      begin
        register_25 <= register_172;
        program_counter <= 16'd75;
      end

      16'd90:
      begin
        register_18 <= 16'd0;
        program_counter <= register_17;
      end

      16'd91:
      begin
        register_31 <= 16'd521;
      end

      16'd92:
      begin
        register_9 <= register_31;
        program_counter <= 16'd2;
        register_7 <= 16'd93;
      end

      16'd93:
      begin
        register_172 <= register_8;
        register_32 <= 16'd0;
        register_33 <= 16'd0;
        register_34 <= 16'd0;
      end

      16'd94:
      begin
        register_172 <= input_eth_rx;
        program_counter <= 94;
        s_input_eth_rx_ack <= 1'b1;
       if (s_input_eth_rx_ack == 1'b1 && input_eth_rx_stb == 1'b1) begin
          s_input_eth_rx_ack <= 1'b0;
          program_counter <= 16'd95;
        end
      end

      16'd95:
      begin
        register_32 <= register_172;
        register_35 <= 16'd530;
      end

      16'd96:
      begin
        register_9 <= register_35;
        program_counter <= 16'd2;
        register_7 <= 16'd97;
      end

      16'd97:
      begin
        register_172 <= register_8;
        register_16 <= register_32;
        program_counter <= 16'd30;
        register_14 <= 16'd98;
      end

      16'd98:
      begin
        register_172 <= register_15;
        register_36 <= 16'd546;
      end

      16'd99:
      begin
        register_9 <= register_36;
        program_counter <= 16'd2;
        register_7 <= 16'd100;
      end

      16'd100:
      begin
        register_172 <= register_8;
      end

      16'd101:
      begin
        register_172 <= 16'd0;
      end

      16'd102:
      begin
        register_33 <= register_172;
        register_172 <= 16'd0;
      end

      16'd103:
      begin
        register_34 <= register_172;
      end

      16'd104:
      begin
        register_172 <= register_34;
        register_173 <= register_32;
      end

      16'd105:
      begin
        register_172 <= $signed(register_172) < $signed(register_173);
      end

      16'd106:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 116;
      end

      16'd107:
      begin
        register_172 <= input_eth_rx;
        program_counter <= 107;
        s_input_eth_rx_ack <= 1'b1;
       if (s_input_eth_rx_ack == 1'b1 && input_eth_rx_stb == 1'b1) begin
          s_input_eth_rx_ack <= 1'b0;
          program_counter <= 16'd108;
        end
      end

      16'd108:
      begin
        register_173 <= register_33;
      end

      16'd109:
      begin
        register_173 <= $signed(register_173) + $signed(register_30);
      end

      16'd110:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_33;
      end

      16'd111:
      begin
        register_172 <= $signed(register_172) + $signed(16'd1);
      end

      16'd112:
      begin
        register_33 <= register_172;
      end

      16'd113:
      begin
        register_172 <= register_34;
      end

      16'd114:
      begin
        register_172 <= $signed(register_172) + $signed(16'd2);
      end

      16'd115:
      begin
        register_34 <= register_172;
        program_counter <= 16'd104;
      end

      16'd116:
      begin
        register_37 <= 16'd548;
      end

      16'd117:
      begin
        register_9 <= register_37;
        program_counter <= 16'd2;
        register_7 <= 16'd118;
      end

      16'd118:
      begin
        register_172 <= register_8;
        register_16 <= 16'd0;
      end

      16'd119:
      begin
        register_16 <= $signed(register_16) + $signed(register_30);
      end

      16'd120:
      begin
        address <= register_16;
      end

      16'd121:
      begin
        register_16 <= data_out;
      end

      16'd122:
      begin
        register_16 <= data_out;
        program_counter <= 16'd30;
        register_14 <= 16'd123;
      end

      16'd123:
      begin
        register_172 <= register_15;
        register_38 <= 16'd554;
      end

      16'd124:
      begin
        register_9 <= register_38;
        program_counter <= 16'd2;
        register_7 <= 16'd125;
      end

      16'd125:
      begin
        register_172 <= register_8;
        register_173 <= register_0;
      end

      16'd126:
      begin
        register_172 <= 16'd0;
      end

      16'd127:
      begin
        register_172 <= $signed(register_172) + $signed(register_30);
      end

      16'd128:
      begin
        address <= register_172;
      end

      16'd129:
      begin
        register_172 <= data_out;
      end

      16'd130:
      begin
        register_172 <= data_out;
      end

      16'd131:
      begin
        register_172 <= $signed(register_172) != $signed(register_173);
      end

      16'd132:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 139;
      end

      16'd133:
      begin
        register_172 <= 16'd0;
      end

      16'd134:
      begin
        register_172 <= $signed(register_172) + $signed(register_30);
      end

      16'd135:
      begin
        address <= register_172;
      end

      16'd136:
      begin
        register_172 <= data_out;
      end

      16'd137:
      begin
        register_172 <= data_out;
      end

      16'd138:
      begin
        register_172 <= $signed(register_172) != $signed(16'd65535);
      end

      16'd139:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 142;
      end

      16'd140:
      begin
        program_counter <= 16'd94;
      end

      16'd141:
      begin
        program_counter <= 16'd142;
      end

      16'd142:
      begin
        register_16 <= 16'd1;
      end

      16'd143:
      begin
        register_16 <= $signed(register_16) + $signed(register_30);
      end

      16'd144:
      begin
        address <= register_16;
      end

      16'd145:
      begin
        register_16 <= data_out;
      end

      16'd146:
      begin
        register_16 <= data_out;
        program_counter <= 16'd30;
        register_14 <= 16'd147;
      end

      16'd147:
      begin
        register_172 <= register_15;
        register_39 <= 16'd556;
      end

      16'd148:
      begin
        register_9 <= register_39;
        program_counter <= 16'd2;
        register_7 <= 16'd149;
      end

      16'd149:
      begin
        register_172 <= register_8;
        register_173 <= register_1;
      end

      16'd150:
      begin
        register_172 <= 16'd1;
      end

      16'd151:
      begin
        register_172 <= $signed(register_172) + $signed(register_30);
      end

      16'd152:
      begin
        address <= register_172;
      end

      16'd153:
      begin
        register_172 <= data_out;
      end

      16'd154:
      begin
        register_172 <= data_out;
      end

      16'd155:
      begin
        register_172 <= $signed(register_172) != $signed(register_173);
      end

      16'd156:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 163;
      end

      16'd157:
      begin
        register_172 <= 16'd1;
      end

      16'd158:
      begin
        register_172 <= $signed(register_172) + $signed(register_30);
      end

      16'd159:
      begin
        address <= register_172;
      end

      16'd160:
      begin
        register_172 <= data_out;
      end

      16'd161:
      begin
        register_172 <= data_out;
      end

      16'd162:
      begin
        register_172 <= $signed(register_172) != $signed(16'd65535);
      end

      16'd163:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 166;
      end

      16'd164:
      begin
        program_counter <= 16'd94;
      end

      16'd165:
      begin
        program_counter <= 16'd166;
      end

      16'd166:
      begin
        register_16 <= 16'd2;
      end

      16'd167:
      begin
        register_16 <= $signed(register_16) + $signed(register_30);
      end

      16'd168:
      begin
        address <= register_16;
      end

      16'd169:
      begin
        register_16 <= data_out;
      end

      16'd170:
      begin
        register_16 <= data_out;
        program_counter <= 16'd30;
        register_14 <= 16'd171;
      end

      16'd171:
      begin
        register_172 <= register_15;
        register_40 <= 16'd558;
      end

      16'd172:
      begin
        register_9 <= register_40;
        program_counter <= 16'd2;
        register_7 <= 16'd173;
      end

      16'd173:
      begin
        register_172 <= register_8;
        register_173 <= register_2;
      end

      16'd174:
      begin
        register_172 <= 16'd2;
      end

      16'd175:
      begin
        register_172 <= $signed(register_172) + $signed(register_30);
      end

      16'd176:
      begin
        address <= register_172;
      end

      16'd177:
      begin
        register_172 <= data_out;
      end

      16'd178:
      begin
        register_172 <= data_out;
      end

      16'd179:
      begin
        register_172 <= $signed(register_172) != $signed(register_173);
      end

      16'd180:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 187;
      end

      16'd181:
      begin
        register_172 <= 16'd2;
      end

      16'd182:
      begin
        register_172 <= $signed(register_172) + $signed(register_30);
      end

      16'd183:
      begin
        address <= register_172;
      end

      16'd184:
      begin
        register_172 <= data_out;
      end

      16'd185:
      begin
        register_172 <= data_out;
      end

      16'd186:
      begin
        register_172 <= $signed(register_172) != $signed(16'd65535);
      end

      16'd187:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 190;
      end

      16'd188:
      begin
        program_counter <= 16'd94;
      end

      16'd189:
      begin
        program_counter <= 16'd190;
      end

      16'd190:
      begin
        register_41 <= 16'd560;
      end

      16'd191:
      begin
        register_9 <= register_41;
        program_counter <= 16'd2;
        register_7 <= 16'd192;
      end

      16'd192:
      begin
        register_172 <= register_8;
      end

      16'd193:
      begin
        register_172 <= 16'd6;
      end

      16'd194:
      begin
        register_172 <= $signed(register_172) + $signed(register_30);
      end

      16'd195:
      begin
        address <= register_172;
      end

      16'd196:
      begin
        register_172 <= data_out;
      end

      16'd197:
      begin
        register_172 <= data_out;
      end

      16'd198:
      begin
        register_172 <= $signed(register_172) == $signed(16'd2054);
      end

      16'd199:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 266;
      end

      16'd200:
      begin
        register_42 <= 16'd570;
      end

      16'd201:
      begin
        register_9 <= register_42;
        program_counter <= 16'd2;
        register_7 <= 16'd202;
      end

      16'd202:
      begin
        register_172 <= register_8;
      end

      16'd203:
      begin
        register_172 <= 16'd10;
      end

      16'd204:
      begin
        register_172 <= $signed(register_172) + $signed(register_30);
      end

      16'd205:
      begin
        address <= register_172;
      end

      16'd206:
      begin
        register_172 <= data_out;
      end

      16'd207:
      begin
        register_172 <= data_out;
      end

      16'd208:
      begin
        register_172 <= $signed(register_172) == $signed(16'd1);
      end

      16'd209:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 264;
      end

      16'd210:
      begin
        register_172 <= 16'd1;
        register_173 <= 16'd7;
        register_19 <= register_6;
        register_20 <= 16'd64;
        register_21 <= 16'd11;
        register_22 <= 16'd12;
        register_23 <= 16'd13;
        register_24 <= 16'd2054;
      end

      16'd211:
      begin
        register_173 <= $signed(register_173) + $signed(register_6);
        register_21 <= $signed(register_21) + $signed(register_30);
        register_22 <= $signed(register_22) + $signed(register_30);
        register_23 <= $signed(register_23) + $signed(register_30);
      end

      16'd212:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= 16'd2048;
        register_173 <= 16'd8;
      end

      16'd213:
      begin
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd214:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= 16'd1540;
        register_173 <= 16'd9;
      end

      16'd215:
      begin
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd216:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= 16'd2;
        register_173 <= 16'd10;
      end

      16'd217:
      begin
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd218:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_0;
        register_173 <= 16'd11;
      end

      16'd219:
      begin
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd220:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_1;
        register_173 <= 16'd12;
      end

      16'd221:
      begin
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd222:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_2;
        register_173 <= 16'd13;
      end

      16'd223:
      begin
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd224:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_3;
        register_173 <= 16'd14;
      end

      16'd225:
      begin
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd226:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_4;
        register_173 <= 16'd15;
      end

      16'd227:
      begin
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd228:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= 16'd11;
        register_173 <= 16'd16;
      end

      16'd229:
      begin
        register_172 <= $signed(register_172) + $signed(register_30);
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd230:
      begin
        address <= register_172;
      end

      16'd231:
      begin
        register_172 <= data_out;
      end

      16'd232:
      begin
        register_172 <= data_out;
      end

      16'd233:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= 16'd12;
        register_173 <= 16'd17;
      end

      16'd234:
      begin
        register_172 <= $signed(register_172) + $signed(register_30);
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd235:
      begin
        address <= register_172;
      end

      16'd236:
      begin
        register_172 <= data_out;
      end

      16'd237:
      begin
        register_172 <= data_out;
      end

      16'd238:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= 16'd13;
        register_173 <= 16'd18;
      end

      16'd239:
      begin
        register_172 <= $signed(register_172) + $signed(register_30);
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd240:
      begin
        address <= register_172;
      end

      16'd241:
      begin
        register_172 <= data_out;
      end

      16'd242:
      begin
        register_172 <= data_out;
      end

      16'd243:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= 16'd14;
        register_173 <= 16'd19;
      end

      16'd244:
      begin
        register_172 <= $signed(register_172) + $signed(register_30);
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd245:
      begin
        address <= register_172;
      end

      16'd246:
      begin
        register_172 <= data_out;
      end

      16'd247:
      begin
        register_172 <= data_out;
      end

      16'd248:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= 16'd15;
        register_173 <= 16'd20;
      end

      16'd249:
      begin
        register_172 <= $signed(register_172) + $signed(register_30);
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd250:
      begin
        address <= register_172;
      end

      16'd251:
      begin
        register_172 <= data_out;
      end

      16'd252:
      begin
        register_172 <= data_out;
      end

      16'd253:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
      end

      16'd254:
      begin
        address <= register_21;
      end

      16'd255:
      begin
        register_21 <= data_out;
      end

      16'd256:
      begin
        register_21 <= data_out;
      end

      16'd257:
      begin
        address <= register_22;
      end

      16'd258:
      begin
        register_22 <= data_out;
      end

      16'd259:
      begin
        register_22 <= data_out;
      end

      16'd260:
      begin
        address <= register_23;
      end

      16'd261:
      begin
        register_23 <= data_out;
      end

      16'd262:
      begin
        register_23 <= data_out;
        program_counter <= 16'd54;
        register_17 <= 16'd263;
      end

      16'd263:
      begin
        register_172 <= register_18;
        program_counter <= 16'd264;
      end

      16'd264:
      begin
        program_counter <= 16'd94;
      end

      16'd265:
      begin
        program_counter <= 16'd266;
      end

      16'd266:
      begin
        program_counter <= 16'd268;
      end

      16'd267:
      begin
        program_counter <= 16'd94;
      end

      16'd268:
      begin
        register_29 <= register_32;
        program_counter <= register_28;
      end

      16'd269:
      begin
        register_53 <= 16'd0;
        register_54 <= 16'd0;
        register_55 <= 16'd655;
        register_56 <= 16'd0;
        register_172 <= 16'd0;
      end

      16'd270:
      begin
        register_56 <= register_172;
      end

      16'd271:
      begin
        register_172 <= register_56;
      end

      16'd272:
      begin
        register_172 <= $signed(register_172) < $signed(16'd16);
      end

      16'd273:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 295;
      end

      16'd274:
      begin
        register_172 <= register_56;
        register_173 <= register_51;
      end

      16'd275:
      begin
        register_172 <= $signed(register_172) + $signed(register_43);
      end

      16'd276:
      begin
        address <= register_172;
      end

      16'd277:
      begin
        register_172 <= data_out;
      end

      16'd278:
      begin
        register_172 <= data_out;
      end

      16'd279:
      begin
        register_172 <= $signed(register_172) == $signed(register_173);
      end

      16'd280:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 287;
      end

      16'd281:
      begin
        register_172 <= register_56;
        register_173 <= register_52;
      end

      16'd282:
      begin
        register_172 <= $signed(register_172) + $signed(register_44);
      end

      16'd283:
      begin
        address <= register_172;
      end

      16'd284:
      begin
        register_172 <= data_out;
      end

      16'd285:
      begin
        register_172 <= data_out;
      end

      16'd286:
      begin
        register_172 <= $signed(register_172) == $signed(register_173);
      end

      16'd287:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 292;
      end

      16'd288:
      begin
        register_57 <= 16'd671;
      end

      16'd289:
      begin
        register_9 <= register_57;
        program_counter <= 16'd2;
        register_7 <= 16'd290;
      end

      16'd290:
      begin
        register_172 <= register_8;
        register_50 <= register_56;
        program_counter <= register_49;
      end

      16'd291:
      begin
        program_counter <= 16'd292;
      end

      16'd292:
      begin
        register_172 <= register_56;
      end

      16'd293:
      begin
        register_172 <= $signed(register_172) + $signed(16'd1);
      end

      16'd294:
      begin
        register_56 <= register_172;
        program_counter <= 16'd271;
      end

      16'd295:
      begin
        register_58 <= 16'd682;
      end

      16'd296:
      begin
        register_9 <= register_58;
        program_counter <= 16'd2;
        register_7 <= 16'd297;
      end

      16'd297:
      begin
        register_172 <= register_8;
        register_173 <= 16'd7;
        register_19 <= register_6;
        register_20 <= 16'd64;
        register_21 <= 16'd65535;
        register_22 <= 16'd65535;
        register_23 <= 16'd65535;
        register_24 <= 16'd2054;
      end

      16'd298:
      begin
        register_172 <= 16'd1;
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd299:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= 16'd2048;
        register_173 <= 16'd8;
      end

      16'd300:
      begin
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd301:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= 16'd1540;
        register_173 <= 16'd9;
      end

      16'd302:
      begin
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd303:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= 16'd1;
        register_173 <= 16'd10;
      end

      16'd304:
      begin
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd305:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_0;
        register_173 <= 16'd11;
      end

      16'd306:
      begin
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd307:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_1;
        register_173 <= 16'd12;
      end

      16'd308:
      begin
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd309:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_2;
        register_173 <= 16'd13;
      end

      16'd310:
      begin
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd311:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_3;
        register_173 <= 16'd14;
      end

      16'd312:
      begin
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd313:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_4;
        register_173 <= 16'd15;
      end

      16'd314:
      begin
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd315:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_51;
        register_173 <= 16'd19;
      end

      16'd316:
      begin
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd317:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_52;
        register_173 <= 16'd20;
      end

      16'd318:
      begin
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd319:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        program_counter <= 16'd54;
        register_17 <= 16'd320;
      end

      16'd320:
      begin
        register_172 <= register_18;
        register_59 <= 16'd694;
      end

      16'd321:
      begin
        register_9 <= register_59;
        program_counter <= 16'd2;
        register_7 <= 16'd322;
      end

      16'd322:
      begin
        register_172 <= register_8;
      end

      16'd323:
      begin
        register_172 <= input_eth_rx;
        program_counter <= 323;
        s_input_eth_rx_ack <= 1'b1;
       if (s_input_eth_rx_ack == 1'b1 && input_eth_rx_stb == 1'b1) begin
          s_input_eth_rx_ack <= 1'b0;
          program_counter <= 16'd324;
        end
      end

      16'd324:
      begin
        register_53 <= register_172;
        register_172 <= 16'd0;
      end

      16'd325:
      begin
        register_56 <= register_172;
        register_172 <= 16'd0;
      end

      16'd326:
      begin
        register_54 <= register_172;
      end

      16'd327:
      begin
        register_172 <= register_54;
        register_173 <= register_53;
      end

      16'd328:
      begin
        register_172 <= $signed(register_172) < $signed(register_173);
      end

      16'd329:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 344;
      end

      16'd330:
      begin
        register_172 <= register_56;
      end

      16'd331:
      begin
        register_172 <= $signed(register_172) < $signed(16'd16);
      end

      16'd332:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 337;
      end

      16'd333:
      begin
        register_172 <= input_eth_rx;
        program_counter <= 333;
        s_input_eth_rx_ack <= 1'b1;
       if (s_input_eth_rx_ack == 1'b1 && input_eth_rx_stb == 1'b1) begin
          s_input_eth_rx_ack <= 1'b0;
          program_counter <= 16'd334;
        end
      end

      16'd334:
      begin
        register_173 <= register_56;
      end

      16'd335:
      begin
        register_173 <= $signed(register_173) + $signed(register_55);
      end

      16'd336:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        program_counter <= 16'd338;
      end

      16'd337:
      begin
        register_172 <= input_eth_rx;
        program_counter <= 337;
        s_input_eth_rx_ack <= 1'b1;
       if (s_input_eth_rx_ack == 1'b1 && input_eth_rx_stb == 1'b1) begin
          s_input_eth_rx_ack <= 1'b0;
          program_counter <= 16'd338;
        end
      end

      16'd338:
      begin
        register_172 <= register_56;
      end

      16'd339:
      begin
        register_172 <= $signed(register_172) + $signed(16'd1);
      end

      16'd340:
      begin
        register_56 <= register_172;
      end

      16'd341:
      begin
        register_172 <= register_54;
      end

      16'd342:
      begin
        register_172 <= $signed(register_172) + $signed(16'd2);
      end

      16'd343:
      begin
        register_54 <= register_172;
        program_counter <= 16'd327;
      end

      16'd344:
      begin
        register_60 <= 16'd707;
      end

      16'd345:
      begin
        register_9 <= register_60;
        program_counter <= 16'd2;
        register_7 <= 16'd346;
      end

      16'd346:
      begin
        register_172 <= register_8;
      end

      16'd347:
      begin
        register_172 <= 16'd6;
      end

      16'd348:
      begin
        register_172 <= $signed(register_172) + $signed(register_55);
      end

      16'd349:
      begin
        address <= register_172;
      end

      16'd350:
      begin
        register_172 <= data_out;
      end

      16'd351:
      begin
        register_172 <= data_out;
      end

      16'd352:
      begin
        register_172 <= $signed(register_172) == $signed(16'd2054);
      end

      16'd353:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 360;
      end

      16'd354:
      begin
        register_172 <= 16'd10;
      end

      16'd355:
      begin
        register_172 <= $signed(register_172) + $signed(register_55);
      end

      16'd356:
      begin
        address <= register_172;
      end

      16'd357:
      begin
        register_172 <= data_out;
      end

      16'd358:
      begin
        register_172 <= data_out;
      end

      16'd359:
      begin
        register_172 <= $signed(register_172) == $signed(16'd2);
      end

      16'd360:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 411;
      end

      16'd361:
      begin
        register_61 <= 16'd719;
      end

      16'd362:
      begin
        register_9 <= register_61;
        program_counter <= 16'd2;
        register_7 <= 16'd363;
      end

      16'd363:
      begin
        register_172 <= register_8;
        register_173 <= register_51;
      end

      16'd364:
      begin
        register_172 <= 16'd14;
      end

      16'd365:
      begin
        register_172 <= $signed(register_172) + $signed(register_55);
      end

      16'd366:
      begin
        address <= register_172;
      end

      16'd367:
      begin
        register_172 <= data_out;
      end

      16'd368:
      begin
        register_172 <= data_out;
      end

      16'd369:
      begin
        register_172 <= $signed(register_172) == $signed(register_173);
      end

      16'd370:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 377;
      end

      16'd371:
      begin
        register_172 <= 16'd15;
        register_173 <= register_52;
      end

      16'd372:
      begin
        register_172 <= $signed(register_172) + $signed(register_55);
      end

      16'd373:
      begin
        address <= register_172;
      end

      16'd374:
      begin
        register_172 <= data_out;
      end

      16'd375:
      begin
        register_172 <= data_out;
      end

      16'd376:
      begin
        register_172 <= $signed(register_172) == $signed(register_173);
      end

      16'd377:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 410;
      end

      16'd378:
      begin
        register_62 <= 16'd733;
      end

      16'd379:
      begin
        register_9 <= register_62;
        program_counter <= 16'd2;
        register_7 <= 16'd380;
      end

      16'd380:
      begin
        register_172 <= register_8;
        register_173 <= register_48;
      end

      16'd381:
      begin
        register_172 <= register_51;
        register_173 <= $signed(register_173) + $signed(register_43);
      end

      16'd382:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_52;
        register_173 <= register_48;
      end

      16'd383:
      begin
        register_173 <= $signed(register_173) + $signed(register_44);
      end

      16'd384:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= 16'd11;
        register_173 <= register_48;
      end

      16'd385:
      begin
        register_172 <= $signed(register_172) + $signed(register_55);
        register_173 <= $signed(register_173) + $signed(register_45);
      end

      16'd386:
      begin
        address <= register_172;
      end

      16'd387:
      begin
        register_172 <= data_out;
      end

      16'd388:
      begin
        register_172 <= data_out;
      end

      16'd389:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= 16'd12;
        register_173 <= register_48;
      end

      16'd390:
      begin
        register_172 <= $signed(register_172) + $signed(register_55);
        register_173 <= $signed(register_173) + $signed(register_46);
      end

      16'd391:
      begin
        address <= register_172;
      end

      16'd392:
      begin
        register_172 <= data_out;
      end

      16'd393:
      begin
        register_172 <= data_out;
      end

      16'd394:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= 16'd13;
        register_173 <= register_48;
      end

      16'd395:
      begin
        register_172 <= $signed(register_172) + $signed(register_55);
        register_173 <= $signed(register_173) + $signed(register_47);
      end

      16'd396:
      begin
        address <= register_172;
      end

      16'd397:
      begin
        register_172 <= data_out;
      end

      16'd398:
      begin
        register_172 <= data_out;
      end

      16'd399:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_48;
      end

      16'd400:
      begin
        register_56 <= register_172;
        register_172 <= register_48;
      end

      16'd401:
      begin
        register_172 <= $signed(register_172) + $signed(16'd1);
      end

      16'd402:
      begin
        register_48 <= register_172;
      end

      16'd403:
      begin
        register_172 <= register_48;
      end

      16'd404:
      begin
        register_172 <= $signed(register_172) == $signed(16'd16);
      end

      16'd405:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 408;
      end

      16'd406:
      begin
        register_172 <= 16'd0;
      end

      16'd407:
      begin
        register_48 <= register_172;
        program_counter <= 16'd408;
      end

      16'd408:
      begin
        register_50 <= register_56;
        program_counter <= register_49;
      end

      16'd409:
      begin
        program_counter <= 16'd410;
      end

      16'd410:
      begin
        program_counter <= 16'd411;
      end

      16'd411:
      begin
        program_counter <= 16'd323;
      end

      16'd412:
      begin
        register_70 <= 16'd749;
      end

      16'd413:
      begin
        register_9 <= register_70;
        program_counter <= 16'd2;
        register_7 <= 16'd414;
      end

      16'd414:
      begin
        register_172 <= register_8;
        register_71 <= 16'd0;
        register_72 <= 16'd0;
        register_73 <= 16'd0;
        register_51 <= register_68;
        register_52 <= register_69;
        program_counter <= 16'd269;
        register_49 <= 16'd415;
      end

      16'd415:
      begin
        register_172 <= register_50;
        register_173 <= 16'd7;
      end

      16'd416:
      begin
        register_73 <= register_172;
        register_172 <= 16'd17664;
        register_173 <= $signed(register_173) + $signed(register_65);
      end

      16'd417:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_66;
        register_173 <= 16'd8;
      end

      16'd418:
      begin
        register_173 <= $signed(register_173) + $signed(register_65);
      end

      16'd419:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= 16'd0;
        register_173 <= 16'd9;
      end

      16'd420:
      begin
        register_173 <= $signed(register_173) + $signed(register_65);
      end

      16'd421:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= 16'd16384;
        register_173 <= 16'd10;
      end

      16'd422:
      begin
        register_173 <= $signed(register_173) + $signed(register_65);
      end

      16'd423:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_67;
        register_173 <= 16'd11;
      end

      16'd424:
      begin
        register_172 <= $signed(16'd65280) | $signed(register_172);
        register_173 <= $signed(register_173) + $signed(register_65);
      end

      16'd425:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= 16'd0;
        register_173 <= 16'd12;
      end

      16'd426:
      begin
        register_173 <= $signed(register_173) + $signed(register_65);
      end

      16'd427:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_3;
        register_173 <= 16'd13;
      end

      16'd428:
      begin
        register_173 <= $signed(register_173) + $signed(register_65);
      end

      16'd429:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_4;
        register_173 <= 16'd14;
      end

      16'd430:
      begin
        register_173 <= $signed(register_173) + $signed(register_65);
      end

      16'd431:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_68;
        register_173 <= 16'd15;
      end

      16'd432:
      begin
        register_173 <= $signed(register_173) + $signed(register_65);
      end

      16'd433:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_69;
        register_173 <= 16'd16;
      end

      16'd434:
      begin
        register_173 <= $signed(register_173) + $signed(register_65);
      end

      16'd435:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_66;
      end

      16'd436:
      begin
        register_172 <= $signed(register_172) + $signed(16'd14);
      end

      16'd437:
      begin
        register_71 <= register_172;
        register_172 <= 16'd10;
      end

      16'd438:
      begin
        s_output_checksum <= register_172;
        program_counter <= 438;
        s_output_checksum_stb <= 1'b1;
        if (s_output_checksum_stb == 1'b1 && output_checksum_ack == 1'b1) begin
          s_output_checksum_stb <= 1'b0;
          program_counter <= 439;
        end
      end

      16'd439:
      begin
        register_172 <= 16'd7;
      end

      16'd440:
      begin
        register_72 <= register_172;
      end

      16'd441:
      begin
        register_172 <= register_72;
      end

      16'd442:
      begin
        register_172 <= $signed(register_172) <= $signed(16'd16);
      end

      16'd443:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 453;
      end

      16'd444:
      begin
        register_172 <= register_72;
      end

      16'd445:
      begin
        register_172 <= $signed(register_172) + $signed(register_65);
      end

      16'd446:
      begin
        address <= register_172;
      end

      16'd447:
      begin
        register_172 <= data_out;
      end

      16'd448:
      begin
        register_172 <= data_out;
      end

      16'd449:
      begin
        s_output_checksum <= register_172;
        program_counter <= 449;
        s_output_checksum_stb <= 1'b1;
        if (s_output_checksum_stb == 1'b1 && output_checksum_ack == 1'b1) begin
          s_output_checksum_stb <= 1'b0;
          program_counter <= 450;
        end
      end

      16'd450:
      begin
        register_172 <= register_72;
      end

      16'd451:
      begin
        register_172 <= $signed(register_172) + $signed(16'd1);
      end

      16'd452:
      begin
        register_72 <= register_172;
        program_counter <= 16'd441;
      end

      16'd453:
      begin
        register_172 <= input_checksum;
        program_counter <= 453;
        s_input_checksum_ack <= 1'b1;
       if (s_input_checksum_ack == 1'b1 && input_checksum_stb == 1'b1) begin
          s_input_checksum_ack <= 1'b0;
          program_counter <= 16'd454;
        end
      end

      16'd454:
      begin
        register_173 <= 16'd12;
      end

      16'd455:
      begin
        register_173 <= $signed(register_173) + $signed(register_65);
      end

      16'd456:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_71;
      end

      16'd457:
      begin
        register_172 <= $signed(register_172) < $signed(16'd64);
      end

      16'd458:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 461;
      end

      16'd459:
      begin
        register_172 <= 16'd64;
      end

      16'd460:
      begin
        register_71 <= register_172;
        program_counter <= 16'd461;
      end

      16'd461:
      begin
        register_19 <= register_65;
        register_20 <= register_71;
        register_21 <= register_73;
        register_22 <= register_73;
        register_23 <= register_73;
        register_24 <= 16'd2048;
      end

      16'd462:
      begin
        register_21 <= $signed(register_21) + $signed(register_45);
        register_22 <= $signed(register_22) + $signed(register_46);
        register_23 <= $signed(register_23) + $signed(register_47);
      end

      16'd463:
      begin
        address <= register_21;
      end

      16'd464:
      begin
        register_21 <= data_out;
      end

      16'd465:
      begin
        register_21 <= data_out;
      end

      16'd466:
      begin
        address <= register_22;
      end

      16'd467:
      begin
        register_22 <= data_out;
      end

      16'd468:
      begin
        register_22 <= data_out;
      end

      16'd469:
      begin
        address <= register_23;
      end

      16'd470:
      begin
        register_23 <= data_out;
      end

      16'd471:
      begin
        register_23 <= data_out;
        program_counter <= 16'd54;
        register_17 <= 16'd472;
      end

      16'd472:
      begin
        register_172 <= register_18;
        register_64 <= 16'd0;
        program_counter <= register_63;
      end

      16'd473:
      begin
        register_77 <= 16'd0;
        register_78 <= 16'd0;
        register_79 <= 16'd0;
        register_80 <= 16'd0;
        register_81 <= 16'd0;
        register_82 <= 16'd0;
        register_83 <= 16'd0;
        register_84 <= 16'd0;
        register_85 <= 16'd0;
        register_86 <= 16'd757;
      end

      16'd474:
      begin
        register_9 <= register_86;
        program_counter <= 16'd2;
        register_7 <= 16'd475;
      end

      16'd475:
      begin
        register_172 <= register_8;
      end

      16'd476:
      begin
        register_30 <= register_76;
        program_counter <= 16'd91;
        register_28 <= 16'd477;
      end

      16'd477:
      begin
        register_172 <= register_29;
      end

      16'd478:
      begin
        register_71 <= register_172;
        register_172 <= 16'd6;
      end

      16'd479:
      begin
        register_172 <= $signed(register_172) + $signed(register_76);
      end

      16'd480:
      begin
        address <= register_172;
      end

      16'd481:
      begin
        register_172 <= data_out;
      end

      16'd482:
      begin
        register_172 <= data_out;
      end

      16'd483:
      begin
        register_172 <= $signed(register_172) == $signed(16'd2048);
      end

      16'd484:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 609;
      end

      16'd485:
      begin
        register_87 <= 16'd765;
      end

      16'd486:
      begin
        register_9 <= register_87;
        program_counter <= 16'd2;
        register_7 <= 16'd487;
      end

      16'd487:
      begin
        register_172 <= register_8;
        register_173 <= register_3;
      end

      16'd488:
      begin
        register_172 <= 16'd15;
      end

      16'd489:
      begin
        register_172 <= $signed(register_172) + $signed(register_76);
      end

      16'd490:
      begin
        address <= register_172;
      end

      16'd491:
      begin
        register_172 <= data_out;
      end

      16'd492:
      begin
        register_172 <= data_out;
      end

      16'd493:
      begin
        register_172 <= $signed(register_172) != $signed(register_173);
      end

      16'd494:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 497;
      end

      16'd495:
      begin
        program_counter <= 16'd476;
      end

      16'd496:
      begin
        program_counter <= 16'd497;
      end

      16'd497:
      begin
        register_172 <= 16'd16;
        register_173 <= register_4;
      end

      16'd498:
      begin
        register_172 <= $signed(register_172) + $signed(register_76);
      end

      16'd499:
      begin
        address <= register_172;
      end

      16'd500:
      begin
        register_172 <= data_out;
      end

      16'd501:
      begin
        register_172 <= data_out;
      end

      16'd502:
      begin
        register_172 <= $signed(register_172) != $signed(register_173);
      end

      16'd503:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 506;
      end

      16'd504:
      begin
        program_counter <= 16'd476;
      end

      16'd505:
      begin
        program_counter <= 16'd506;
      end

      16'd506:
      begin
        register_88 <= 16'd769;
      end

      16'd507:
      begin
        register_9 <= register_88;
        program_counter <= 16'd2;
        register_7 <= 16'd508;
      end

      16'd508:
      begin
        register_172 <= register_8;
      end

      16'd509:
      begin
        register_172 <= 16'd11;
      end

      16'd510:
      begin
        register_172 <= $signed(register_172) + $signed(register_76);
      end

      16'd511:
      begin
        address <= register_172;
      end

      16'd512:
      begin
        register_172 <= data_out;
      end

      16'd513:
      begin
        register_172 <= data_out;
      end

      16'd514:
      begin
        register_172 <= $signed(register_172) & $signed(16'd255);
      end

      16'd515:
      begin
        register_172 <= $signed(register_172) == $signed(16'd1);
      end

      16'd516:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 598;
      end

      16'd517:
      begin
        register_172 <= 16'd7;
        register_89 <= 16'd786;
      end

      16'd518:
      begin
        register_172 <= $signed(register_172) + $signed(register_76);
        register_9 <= register_89;
      end

      16'd519:
      begin
        address <= register_172;
      end

      16'd520:
      begin
        register_172 <= data_out;
      end

      16'd521:
      begin
        register_172 <= data_out;
      end

      16'd522:
      begin
        register_172 <= $signed(register_172) >>> $signed(16'd8);
      end

      16'd523:
      begin
        register_172 <= $signed(register_172) & $signed(16'd15);
      end

      16'd524:
      begin
        register_172 <= $signed(register_172) << $signed(16'd1);
      end

      16'd525:
      begin
        register_79 <= register_172;
      end

      16'd526:
      begin
        register_172 <= register_79;
        register_173 <= register_79;
      end

      16'd527:
      begin
        register_172 <= $signed(register_172) + $signed(16'd7);
      end

      16'd528:
      begin
        register_80 <= register_172;
        register_172 <= 16'd8;
      end

      16'd529:
      begin
        register_172 <= $signed(register_172) + $signed(register_76);
      end

      16'd530:
      begin
        address <= register_172;
      end

      16'd531:
      begin
        register_172 <= data_out;
      end

      16'd532:
      begin
        register_172 <= data_out;
      end

      16'd533:
      begin
        register_78 <= register_172;
      end

      16'd534:
      begin
        register_172 <= register_78;
      end

      16'd535:
      begin
        register_172 <= $signed(register_172) + $signed(16'd1);
      end

      16'd536:
      begin
        register_172 <= $signed(register_172) >>> $signed(16'd1);
      end

      16'd537:
      begin
        register_172 <= $signed(register_172) - $signed(register_173);
      end

      16'd538:
      begin
        register_81 <= register_172;
        register_172 <= register_80;
      end

      16'd539:
      begin
        register_173 <= register_81;
      end

      16'd540:
      begin
        register_172 <= $signed(register_172) + $signed(register_173);
      end

      16'd541:
      begin
        register_172 <= $signed(register_172) - $signed(16'd1);
      end

      16'd542:
      begin
        register_85 <= register_172;
        program_counter <= 16'd2;
        register_7 <= 16'd543;
      end

      16'd543:
      begin
        register_172 <= register_8;
      end

      16'd544:
      begin
        register_172 <= register_80;
      end

      16'd545:
      begin
        register_172 <= $signed(register_172) + $signed(register_76);
      end

      16'd546:
      begin
        address <= register_172;
      end

      16'd547:
      begin
        register_172 <= data_out;
      end

      16'd548:
      begin
        register_172 <= data_out;
      end

      16'd549:
      begin
        register_172 <= $signed(register_172) == $signed(16'd2048);
      end

      16'd550:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 597;
      end

      16'd551:
      begin
        register_90 <= 16'd792;
      end

      16'd552:
      begin
        register_9 <= register_90;
        program_counter <= 16'd2;
        register_7 <= 16'd553;
      end

      16'd553:
      begin
        register_172 <= register_8;
      end

      16'd554:
      begin
        register_172 <= 16'd19;
      end

      16'd555:
      begin
        register_84 <= register_172;
        register_172 <= register_81;
      end

      16'd556:
      begin
        s_output_checksum <= register_172;
        program_counter <= 556;
        s_output_checksum_stb <= 1'b1;
        if (s_output_checksum_stb == 1'b1 && output_checksum_ack == 1'b1) begin
          s_output_checksum_stb <= 1'b0;
          program_counter <= 557;
        end
      end

      16'd557:
      begin
        register_172 <= 16'd0;
      end

      16'd558:
      begin
        s_output_checksum <= register_172;
        program_counter <= 558;
        s_output_checksum_stb <= 1'b1;
        if (s_output_checksum_stb == 1'b1 && output_checksum_ack == 1'b1) begin
          s_output_checksum_stb <= 1'b0;
          program_counter <= 559;
        end
      end

      16'd559:
      begin
        register_172 <= 16'd0;
      end

      16'd560:
      begin
        s_output_checksum <= register_172;
        program_counter <= 560;
        s_output_checksum_stb <= 1'b1;
        if (s_output_checksum_stb == 1'b1 && output_checksum_ack == 1'b1) begin
          s_output_checksum_stb <= 1'b0;
          program_counter <= 561;
        end
      end

      16'd561:
      begin
        register_172 <= register_80;
      end

      16'd562:
      begin
        register_172 <= $signed(register_172) + $signed(16'd2);
      end

      16'd563:
      begin
        register_83 <= register_172;
      end

      16'd564:
      begin
        register_172 <= register_83;
        register_173 <= register_85;
      end

      16'd565:
      begin
        register_172 <= $signed(register_172) <= $signed(register_173);
      end

      16'd566:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 583;
      end

      16'd567:
      begin
        register_172 <= register_83;
      end

      16'd568:
      begin
        register_172 <= $signed(register_172) + $signed(register_76);
      end

      16'd569:
      begin
        address <= register_172;
      end

      16'd570:
      begin
        register_172 <= data_out;
      end

      16'd571:
      begin
        register_172 <= data_out;
      end

      16'd572:
      begin
        register_82 <= register_172;
      end

      16'd573:
      begin
        register_172 <= register_82;
      end

      16'd574:
      begin
        s_output_checksum <= register_172;
        program_counter <= 574;
        s_output_checksum_stb <= 1'b1;
        if (s_output_checksum_stb == 1'b1 && output_checksum_ack == 1'b1) begin
          s_output_checksum_stb <= 1'b0;
          program_counter <= 575;
        end
      end

      16'd575:
      begin
        register_172 <= register_82;
        register_173 <= register_84;
      end

      16'd576:
      begin
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd577:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_84;
      end

      16'd578:
      begin
        register_172 <= $signed(register_172) + $signed(16'd1);
      end

      16'd579:
      begin
        register_84 <= register_172;
      end

      16'd580:
      begin
        register_172 <= register_83;
      end

      16'd581:
      begin
        register_172 <= $signed(register_172) + $signed(16'd1);
      end

      16'd582:
      begin
        register_83 <= register_172;
        program_counter <= 16'd564;
      end

      16'd583:
      begin
        register_172 <= 16'd0;
        register_173 <= 16'd17;
      end

      16'd584:
      begin
        register_173 <= $signed(register_173) + $signed(register_6);
      end

      16'd585:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
      end

      16'd586:
      begin
        register_172 <= input_checksum;
        program_counter <= 586;
        s_input_checksum_ack <= 1'b1;
       if (s_input_checksum_ack == 1'b1 && input_checksum_stb == 1'b1) begin
          s_input_checksum_ack <= 1'b0;
          program_counter <= 16'd587;
        end
      end

      16'd587:
      begin
        register_173 <= 16'd18;
        register_65 <= register_6;
        register_66 <= register_78;
        register_67 <= 16'd1;
        register_68 <= 16'd13;
        register_69 <= 16'd14;
      end

      16'd588:
      begin
        register_173 <= $signed(register_173) + $signed(register_6);
        register_68 <= $signed(register_68) + $signed(register_76);
        register_69 <= $signed(register_69) + $signed(register_76);
      end

      16'd589:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
      end

      16'd590:
      begin
        address <= register_68;
      end

      16'd591:
      begin
        register_68 <= data_out;
      end

      16'd592:
      begin
        register_68 <= data_out;
      end

      16'd593:
      begin
        address <= register_69;
      end

      16'd594:
      begin
        register_69 <= data_out;
      end

      16'd595:
      begin
        register_69 <= data_out;
        program_counter <= 16'd412;
        register_63 <= 16'd596;
      end

      16'd596:
      begin
        register_172 <= register_64;
        program_counter <= 16'd597;
      end

      16'd597:
      begin
        program_counter <= 16'd608;
      end

      16'd598:
      begin
        register_172 <= 16'd11;
      end

      16'd599:
      begin
        register_172 <= $signed(register_172) + $signed(register_76);
      end

      16'd600:
      begin
        address <= register_172;
      end

      16'd601:
      begin
        register_172 <= data_out;
      end

      16'd602:
      begin
        register_172 <= data_out;
      end

      16'd603:
      begin
        register_172 <= $signed(register_172) & $signed(16'd255);
      end

      16'd604:
      begin
        register_172 <= $signed(register_172) == $signed(16'd6);
      end

      16'd605:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 608;
      end

      16'd606:
      begin
        register_75 <= register_71;
        program_counter <= register_74;
      end

      16'd607:
      begin
        program_counter <= 16'd608;
      end

      16'd608:
      begin
        program_counter <= 16'd612;
      end

      16'd609:
      begin
        register_91 <= 16'd806;
      end

      16'd610:
      begin
        register_9 <= register_91;
        program_counter <= 16'd2;
        register_7 <= 16'd611;
      end

      16'd611:
      begin
        register_172 <= register_8;
      end

      16'd612:
      begin
        program_counter <= 16'd476;
      end

      16'd613:
      begin
        register_124 <= 16'd812;
      end

      16'd614:
      begin
        register_9 <= register_124;
        program_counter <= 16'd2;
        register_7 <= 16'd615;
      end

      16'd615:
      begin
        register_172 <= register_8;
        register_125 <= 16'd17;
        register_126 <= 16'd0;
        register_127 <= 16'd0;
        register_128 <= 16'd0;
      end

      16'd616:
      begin
        register_172 <= register_94;
        register_173 <= register_125;
      end

      16'd617:
      begin
        register_173 <= $signed(register_173) + $signed(16'd0);
      end

      16'd618:
      begin
        register_173 <= $signed(register_173) + $signed(register_122);
      end

      16'd619:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_95;
        register_173 <= register_125;
      end

      16'd620:
      begin
        register_173 <= $signed(register_173) + $signed(16'd1);
      end

      16'd621:
      begin
        register_173 <= $signed(register_173) + $signed(register_122);
      end

      16'd622:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_96;
        register_173 <= register_125;
      end

      16'd623:
      begin
        register_173 <= $signed(register_173) + $signed(16'd2);
      end

      16'd624:
      begin
        register_173 <= $signed(register_173) + $signed(register_122);
      end

      16'd625:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_97;
        register_173 <= register_125;
      end

      16'd626:
      begin
        register_173 <= $signed(register_173) + $signed(16'd3);
      end

      16'd627:
      begin
        register_173 <= $signed(register_173) + $signed(register_122);
      end

      16'd628:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_98;
        register_173 <= register_125;
      end

      16'd629:
      begin
        register_173 <= $signed(register_173) + $signed(16'd4);
      end

      16'd630:
      begin
        register_173 <= $signed(register_173) + $signed(register_122);
      end

      16'd631:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_99;
        register_173 <= register_125;
      end

      16'd632:
      begin
        register_173 <= $signed(register_173) + $signed(16'd5);
      end

      16'd633:
      begin
        register_173 <= $signed(register_173) + $signed(register_122);
      end

      16'd634:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= 16'd20480;
        register_173 <= register_125;
      end

      16'd635:
      begin
        register_173 <= $signed(register_173) + $signed(16'd6);
      end

      16'd636:
      begin
        register_173 <= $signed(register_173) + $signed(register_122);
      end

      16'd637:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_100;
        register_173 <= register_125;
      end

      16'd638:
      begin
        register_173 <= $signed(register_173) + $signed(16'd7);
      end

      16'd639:
      begin
        register_173 <= $signed(register_173) + $signed(register_122);
      end

      16'd640:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= 16'd0;
        register_173 <= register_125;
      end

      16'd641:
      begin
        register_173 <= $signed(register_173) + $signed(16'd8);
      end

      16'd642:
      begin
        register_173 <= $signed(register_173) + $signed(register_122);
      end

      16'd643:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= 16'd0;
        register_173 <= register_125;
      end

      16'd644:
      begin
        register_173 <= $signed(register_173) + $signed(16'd9);
      end

      16'd645:
      begin
        register_173 <= $signed(register_173) + $signed(register_122);
      end

      16'd646:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        register_172 <= register_101;
      end

      16'd647:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 656;
      end

      16'd648:
      begin
        register_172 <= register_125;
        register_173 <= register_125;
      end

      16'd649:
      begin
        register_172 <= $signed(register_172) + $signed(16'd6);
        register_173 <= $signed(register_173) + $signed(16'd6);
      end

      16'd650:
      begin
        register_172 <= $signed(register_172) + $signed(register_122);
        register_173 <= $signed(register_173) + $signed(register_122);
      end

      16'd651:
      begin
        address <= register_172;
      end

      16'd652:
      begin
        register_172 <= data_out;
      end

      16'd653:
      begin
        register_172 <= data_out;
      end

      16'd654:
      begin
        register_172 <= $signed(register_172) | $signed(16'd1);
      end

      16'd655:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        program_counter <= 16'd656;
      end

      16'd656:
      begin
        register_172 <= register_102;
      end

      16'd657:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 666;
      end

      16'd658:
      begin
        register_172 <= register_125;
        register_173 <= register_125;
      end

      16'd659:
      begin
        register_172 <= $signed(register_172) + $signed(16'd6);
        register_173 <= $signed(register_173) + $signed(16'd6);
      end

      16'd660:
      begin
        register_172 <= $signed(register_172) + $signed(register_122);
        register_173 <= $signed(register_173) + $signed(register_122);
      end

      16'd661:
      begin
        address <= register_172;
      end

      16'd662:
      begin
        register_172 <= data_out;
      end

      16'd663:
      begin
        register_172 <= data_out;
      end

      16'd664:
      begin
        register_172 <= $signed(register_172) | $signed(16'd2);
      end

      16'd665:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        program_counter <= 16'd666;
      end

      16'd666:
      begin
        register_172 <= register_103;
      end

      16'd667:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 676;
      end

      16'd668:
      begin
        register_172 <= register_125;
        register_173 <= register_125;
      end

      16'd669:
      begin
        register_172 <= $signed(register_172) + $signed(16'd6);
        register_173 <= $signed(register_173) + $signed(16'd6);
      end

      16'd670:
      begin
        register_172 <= $signed(register_172) + $signed(register_122);
        register_173 <= $signed(register_173) + $signed(register_122);
      end

      16'd671:
      begin
        address <= register_172;
      end

      16'd672:
      begin
        register_172 <= data_out;
      end

      16'd673:
      begin
        register_172 <= data_out;
      end

      16'd674:
      begin
        register_172 <= $signed(register_172) | $signed(16'd4);
      end

      16'd675:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        program_counter <= 16'd676;
      end

      16'd676:
      begin
        register_172 <= register_104;
      end

      16'd677:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 686;
      end

      16'd678:
      begin
        register_172 <= register_125;
        register_173 <= register_125;
      end

      16'd679:
      begin
        register_172 <= $signed(register_172) + $signed(16'd6);
        register_173 <= $signed(register_173) + $signed(16'd6);
      end

      16'd680:
      begin
        register_172 <= $signed(register_172) + $signed(register_122);
        register_173 <= $signed(register_173) + $signed(register_122);
      end

      16'd681:
      begin
        address <= register_172;
      end

      16'd682:
      begin
        register_172 <= data_out;
      end

      16'd683:
      begin
        register_172 <= data_out;
      end

      16'd684:
      begin
        register_172 <= $signed(register_172) | $signed(16'd8);
      end

      16'd685:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        program_counter <= 16'd686;
      end

      16'd686:
      begin
        register_172 <= register_105;
      end

      16'd687:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 696;
      end

      16'd688:
      begin
        register_172 <= register_125;
        register_173 <= register_125;
      end

      16'd689:
      begin
        register_172 <= $signed(register_172) + $signed(16'd6);
        register_173 <= $signed(register_173) + $signed(16'd6);
      end

      16'd690:
      begin
        register_172 <= $signed(register_172) + $signed(register_122);
        register_173 <= $signed(register_173) + $signed(register_122);
      end

      16'd691:
      begin
        address <= register_172;
      end

      16'd692:
      begin
        register_172 <= data_out;
      end

      16'd693:
      begin
        register_172 <= data_out;
      end

      16'd694:
      begin
        register_172 <= $signed(register_172) | $signed(16'd16);
      end

      16'd695:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        program_counter <= 16'd696;
      end

      16'd696:
      begin
        register_172 <= register_106;
      end

      16'd697:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 706;
      end

      16'd698:
      begin
        register_172 <= register_125;
        register_173 <= register_125;
      end

      16'd699:
      begin
        register_172 <= $signed(register_172) + $signed(16'd6);
        register_173 <= $signed(register_173) + $signed(16'd6);
      end

      16'd700:
      begin
        register_172 <= $signed(register_172) + $signed(register_122);
        register_173 <= $signed(register_173) + $signed(register_122);
      end

      16'd701:
      begin
        address <= register_172;
      end

      16'd702:
      begin
        register_172 <= data_out;
      end

      16'd703:
      begin
        register_172 <= data_out;
      end

      16'd704:
      begin
        register_172 <= $signed(register_172) | $signed(16'd32);
      end

      16'd705:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        program_counter <= 16'd706;
      end

      16'd706:
      begin
        register_172 <= register_123;
      end

      16'd707:
      begin
        register_172 <= $signed(register_172) + $signed(16'd20);
      end

      16'd708:
      begin
        register_172 <= $signed(register_172) + $signed(16'd12);
      end

      16'd709:
      begin
        register_172 <= $signed(register_172) + $signed(16'd1);
      end

      16'd710:
      begin
        register_172 <= $signed(register_172) >>> $signed(16'd1);
      end

      16'd711:
      begin
        register_126 <= register_172;
      end

      16'd712:
      begin
        register_172 <= register_126;
      end

      16'd713:
      begin
        s_output_checksum <= register_172;
        program_counter <= 713;
        s_output_checksum_stb <= 1'b1;
        if (s_output_checksum_stb == 1'b1 && output_checksum_ack == 1'b1) begin
          s_output_checksum_stb <= 1'b0;
          program_counter <= 714;
        end
      end

      16'd714:
      begin
        register_172 <= register_3;
      end

      16'd715:
      begin
        s_output_checksum <= register_172;
        program_counter <= 715;
        s_output_checksum_stb <= 1'b1;
        if (s_output_checksum_stb == 1'b1 && output_checksum_ack == 1'b1) begin
          s_output_checksum_stb <= 1'b0;
          program_counter <= 716;
        end
      end

      16'd716:
      begin
        register_172 <= register_4;
      end

      16'd717:
      begin
        s_output_checksum <= register_172;
        program_counter <= 717;
        s_output_checksum_stb <= 1'b1;
        if (s_output_checksum_stb == 1'b1 && output_checksum_ack == 1'b1) begin
          s_output_checksum_stb <= 1'b0;
          program_counter <= 718;
        end
      end

      16'd718:
      begin
        register_172 <= register_92;
      end

      16'd719:
      begin
        s_output_checksum <= register_172;
        program_counter <= 719;
        s_output_checksum_stb <= 1'b1;
        if (s_output_checksum_stb == 1'b1 && output_checksum_ack == 1'b1) begin
          s_output_checksum_stb <= 1'b0;
          program_counter <= 720;
        end
      end

      16'd720:
      begin
        register_172 <= register_93;
      end

      16'd721:
      begin
        s_output_checksum <= register_172;
        program_counter <= 721;
        s_output_checksum_stb <= 1'b1;
        if (s_output_checksum_stb == 1'b1 && output_checksum_ack == 1'b1) begin
          s_output_checksum_stb <= 1'b0;
          program_counter <= 722;
        end
      end

      16'd722:
      begin
        register_172 <= 16'd6;
      end

      16'd723:
      begin
        s_output_checksum <= register_172;
        program_counter <= 723;
        s_output_checksum_stb <= 1'b1;
        if (s_output_checksum_stb == 1'b1 && output_checksum_ack == 1'b1) begin
          s_output_checksum_stb <= 1'b0;
          program_counter <= 724;
        end
      end

      16'd724:
      begin
        register_172 <= register_123;
      end

      16'd725:
      begin
        register_172 <= $signed(register_172) + $signed(16'd20);
      end

      16'd726:
      begin
        s_output_checksum <= register_172;
        program_counter <= 726;
        s_output_checksum_stb <= 1'b1;
        if (s_output_checksum_stb == 1'b1 && output_checksum_ack == 1'b1) begin
          s_output_checksum_stb <= 1'b0;
          program_counter <= 727;
        end
      end

      16'd727:
      begin
        register_172 <= register_123;
      end

      16'd728:
      begin
        register_172 <= $signed(register_172) + $signed(16'd20);
      end

      16'd729:
      begin
        register_172 <= $signed(register_172) + $signed(16'd1);
      end

      16'd730:
      begin
        register_172 <= $signed(register_172) >>> $signed(16'd1);
      end

      16'd731:
      begin
        register_127 <= register_172;
        register_172 <= register_125;
      end

      16'd732:
      begin
        register_128 <= register_172;
        register_172 <= 16'd0;
      end

      16'd733:
      begin
        register_82 <= register_172;
      end

      16'd734:
      begin
        register_172 <= register_82;
        register_173 <= register_127;
      end

      16'd735:
      begin
        register_172 <= $signed(register_172) < $signed(register_173);
      end

      16'd736:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 749;
      end

      16'd737:
      begin
        register_172 <= register_128;
      end

      16'd738:
      begin
        register_172 <= $signed(register_172) + $signed(register_122);
      end

      16'd739:
      begin
        address <= register_172;
      end

      16'd740:
      begin
        register_172 <= data_out;
      end

      16'd741:
      begin
        register_172 <= data_out;
      end

      16'd742:
      begin
        s_output_checksum <= register_172;
        program_counter <= 742;
        s_output_checksum_stb <= 1'b1;
        if (s_output_checksum_stb == 1'b1 && output_checksum_ack == 1'b1) begin
          s_output_checksum_stb <= 1'b0;
          program_counter <= 743;
        end
      end

      16'd743:
      begin
        register_172 <= register_128;
      end

      16'd744:
      begin
        register_172 <= $signed(register_172) + $signed(16'd1);
      end

      16'd745:
      begin
        register_128 <= register_172;
      end

      16'd746:
      begin
        register_172 <= register_82;
      end

      16'd747:
      begin
        register_172 <= $signed(register_172) + $signed(16'd1);
      end

      16'd748:
      begin
        register_82 <= register_172;
        program_counter <= 16'd734;
      end

      16'd749:
      begin
        register_172 <= input_checksum;
        program_counter <= 749;
        s_input_checksum_ack <= 1'b1;
       if (s_input_checksum_ack == 1'b1 && input_checksum_stb == 1'b1) begin
          s_input_checksum_ack <= 1'b0;
          program_counter <= 16'd750;
        end
      end

      16'd750:
      begin
        register_173 <= register_125;
        register_65 <= register_122;
        register_66 <= register_123;
        register_67 <= 16'd6;
        register_68 <= register_92;
        register_69 <= register_93;
      end

      16'd751:
      begin
        register_173 <= $signed(register_173) + $signed(16'd8);
        register_66 <= $signed(register_66) + $signed(16'd40);
      end

      16'd752:
      begin
        register_173 <= $signed(register_173) + $signed(register_122);
      end

      16'd753:
      begin
        address <= register_173;
        data_in <= register_172;
        write_enable <= 1'b1;
        program_counter <= 16'd412;
        register_63 <= 16'd754;
      end

      16'd754:
      begin
        register_172 <= register_64;
        register_121 <= 16'd0;
        program_counter <= register_120;
      end

      16'd755:
      begin
        register_132 <= 16'd821;
      end

      16'd756:
      begin
        register_9 <= register_132;
        program_counter <= 16'd2;
        register_7 <= 16'd757;
      end

      16'd757:
      begin
        register_172 <= register_8;
        register_133 <= 16'd0;
        register_134 <= 16'd0;
        register_135 <= 16'd0;
        register_136 <= 16'd0;
        register_137 <= 16'd0;
        register_138 <= 16'd0;
        register_139 <= 16'd0;
        register_140 <= 16'd0;
        register_76 <= register_131;
        program_counter <= 16'd473;
        register_74 <= 16'd758;
      end

      16'd758:
      begin
        register_172 <= register_75;
        register_141 <= 16'd830;
      end

      16'd759:
      begin
        register_133 <= register_172;
        register_172 <= 16'd7;
        register_9 <= register_141;
      end

      16'd760:
      begin
        register_172 <= $signed(register_172) + $signed(register_131);
      end

      16'd761:
      begin
        address <= register_172;
      end

      16'd762:
      begin
        register_172 <= data_out;
      end

      16'd763:
      begin
        register_172 <= data_out;
      end

      16'd764:
      begin
        register_172 <= $signed(register_172) >>> $signed(16'd8);
      end

      16'd765:
      begin
        register_172 <= $signed(register_172) & $signed(16'd15);
      end

      16'd766:
      begin
        register_172 <= $signed(register_172) << $signed(16'd1);
      end

      16'd767:
      begin
        register_134 <= register_172;
      end

      16'd768:
      begin
        register_172 <= register_134;
        register_173 <= register_134;
      end

      16'd769:
      begin
        register_172 <= $signed(register_172) + $signed(16'd7);
      end

      16'd770:
      begin
        register_135 <= register_172;
        register_172 <= 16'd8;
      end

      16'd771:
      begin
        register_172 <= $signed(register_172) + $signed(register_131);
      end

      16'd772:
      begin
        address <= register_172;
      end

      16'd773:
      begin
        register_172 <= data_out;
      end

      16'd774:
      begin
        register_172 <= data_out;
      end

      16'd775:
      begin
        register_136 <= register_172;
      end

      16'd776:
      begin
        register_172 <= register_136;
      end

      16'd777:
      begin
        register_172 <= $signed(register_172) + $signed(16'd1);
      end

      16'd778:
      begin
        register_172 <= $signed(register_172) >>> $signed(16'd1);
      end

      16'd779:
      begin
        register_172 <= $signed(register_172) - $signed(register_173);
      end

      16'd780:
      begin
        register_137 <= register_172;
        register_172 <= register_135;
      end

      16'd781:
      begin
        register_173 <= register_137;
      end

      16'd782:
      begin
        register_172 <= $signed(register_172) + $signed(register_173);
      end

      16'd783:
      begin
        register_172 <= $signed(register_172) - $signed(16'd1);
      end

      16'd784:
      begin
        register_138 <= register_172;
        register_172 <= register_135;
      end

      16'd785:
      begin
        register_172 <= $signed(register_172) + $signed(16'd6);
      end

      16'd786:
      begin
        register_172 <= $signed(register_172) + $signed(register_131);
      end

      16'd787:
      begin
        address <= register_172;
      end

      16'd788:
      begin
        register_172 <= data_out;
      end

      16'd789:
      begin
        register_172 <= data_out;
      end

      16'd790:
      begin
        register_172 <= $signed(register_172) & $signed(16'd61440);
      end

      16'd791:
      begin
        register_172 <= $signed(register_172) >>> $signed(16'd11);
      end

      16'd792:
      begin
        register_139 <= register_172;
        register_172 <= register_137;
      end

      16'd793:
      begin
        register_173 <= register_139;
      end

      16'd794:
      begin
        register_172 <= $signed(register_172) - $signed(register_173);
      end

      16'd795:
      begin
        register_140 <= register_172;
        register_172 <= register_135;
      end

      16'd796:
      begin
        register_172 <= $signed(register_172) + $signed(16'd0);
      end

      16'd797:
      begin
        register_172 <= $signed(register_172) + $signed(register_131);
      end

      16'd798:
      begin
        address <= register_172;
      end

      16'd799:
      begin
        register_172 <= data_out;
      end

      16'd800:
      begin
        register_172 <= data_out;
      end

      16'd801:
      begin
        register_107 <= register_172;
        register_172 <= register_135;
      end

      16'd802:
      begin
        register_172 <= $signed(register_172) + $signed(16'd1);
      end

      16'd803:
      begin
        register_172 <= $signed(register_172) + $signed(register_131);
      end

      16'd804:
      begin
        address <= register_172;
      end

      16'd805:
      begin
        register_172 <= data_out;
      end

      16'd806:
      begin
        register_172 <= data_out;
      end

      16'd807:
      begin
        register_108 <= register_172;
        register_172 <= register_135;
      end

      16'd808:
      begin
        register_172 <= $signed(register_172) + $signed(16'd2);
      end

      16'd809:
      begin
        register_172 <= $signed(register_172) + $signed(register_131);
      end

      16'd810:
      begin
        address <= register_172;
      end

      16'd811:
      begin
        register_172 <= data_out;
      end

      16'd812:
      begin
        register_172 <= data_out;
      end

      16'd813:
      begin
        register_109 <= register_172;
        register_172 <= register_135;
      end

      16'd814:
      begin
        register_172 <= $signed(register_172) + $signed(16'd3);
      end

      16'd815:
      begin
        register_172 <= $signed(register_172) + $signed(register_131);
      end

      16'd816:
      begin
        address <= register_172;
      end

      16'd817:
      begin
        register_172 <= data_out;
      end

      16'd818:
      begin
        register_172 <= data_out;
      end

      16'd819:
      begin
        register_110 <= register_172;
        register_172 <= register_135;
      end

      16'd820:
      begin
        register_172 <= $signed(register_172) + $signed(16'd4);
      end

      16'd821:
      begin
        register_172 <= $signed(register_172) + $signed(register_131);
      end

      16'd822:
      begin
        address <= register_172;
      end

      16'd823:
      begin
        register_172 <= data_out;
      end

      16'd824:
      begin
        register_172 <= data_out;
      end

      16'd825:
      begin
        register_111 <= register_172;
        register_172 <= register_135;
      end

      16'd826:
      begin
        register_172 <= $signed(register_172) + $signed(16'd5);
      end

      16'd827:
      begin
        register_172 <= $signed(register_172) + $signed(register_131);
      end

      16'd828:
      begin
        address <= register_172;
      end

      16'd829:
      begin
        register_172 <= data_out;
      end

      16'd830:
      begin
        register_172 <= data_out;
      end

      16'd831:
      begin
        register_112 <= register_172;
        register_172 <= register_135;
      end

      16'd832:
      begin
        register_172 <= $signed(register_172) + $signed(16'd7);
      end

      16'd833:
      begin
        register_172 <= $signed(register_172) + $signed(register_131);
      end

      16'd834:
      begin
        address <= register_172;
      end

      16'd835:
      begin
        register_172 <= data_out;
      end

      16'd836:
      begin
        register_172 <= data_out;
      end

      16'd837:
      begin
        register_113 <= register_172;
        program_counter <= 16'd2;
        register_7 <= 16'd838;
      end

      16'd838:
      begin
        register_172 <= register_8;
        register_16 <= register_107;
        program_counter <= 16'd30;
        register_14 <= 16'd839;
      end

      16'd839:
      begin
        register_172 <= register_15;
        register_142 <= 16'd839;
      end

      16'd840:
      begin
        register_9 <= register_142;
        program_counter <= 16'd2;
        register_7 <= 16'd841;
      end

      16'd841:
      begin
        register_172 <= register_8;
        register_143 <= 16'd841;
      end

      16'd842:
      begin
        register_9 <= register_143;
        program_counter <= 16'd2;
        register_7 <= 16'd843;
      end

      16'd843:
      begin
        register_172 <= register_8;
        register_16 <= register_108;
        program_counter <= 16'd30;
        register_14 <= 16'd844;
      end

      16'd844:
      begin
        register_172 <= register_15;
        register_144 <= 16'd848;
      end

      16'd845:
      begin
        register_9 <= register_144;
        program_counter <= 16'd2;
        register_7 <= 16'd846;
      end

      16'd846:
      begin
        register_172 <= register_8;
        register_145 <= 16'd850;
      end

      16'd847:
      begin
        register_9 <= register_145;
        program_counter <= 16'd2;
        register_7 <= 16'd848;
      end

      16'd848:
      begin
        register_172 <= register_8;
        register_16 <= register_109;
        program_counter <= 16'd30;
        register_14 <= 16'd849;
      end

      16'd849:
      begin
        register_172 <= register_15;
        register_146 <= 16'd859;
      end

      16'd850:
      begin
        register_9 <= register_146;
        program_counter <= 16'd2;
        register_7 <= 16'd851;
      end

      16'd851:
      begin
        register_172 <= register_8;
        register_147 <= 16'd861;
      end

      16'd852:
      begin
        register_9 <= register_147;
        program_counter <= 16'd2;
        register_7 <= 16'd853;
      end

      16'd853:
      begin
        register_172 <= register_8;
        register_16 <= register_110;
        program_counter <= 16'd30;
        register_14 <= 16'd854;
      end

      16'd854:
      begin
        register_172 <= register_15;
        register_148 <= 16'd870;
      end

      16'd855:
      begin
        register_9 <= register_148;
        program_counter <= 16'd2;
        register_7 <= 16'd856;
      end

      16'd856:
      begin
        register_172 <= register_8;
        register_149 <= 16'd872;
      end

      16'd857:
      begin
        register_9 <= register_149;
        program_counter <= 16'd2;
        register_7 <= 16'd858;
      end

      16'd858:
      begin
        register_172 <= register_8;
        register_16 <= register_111;
        program_counter <= 16'd30;
        register_14 <= 16'd859;
      end

      16'd859:
      begin
        register_172 <= register_15;
        register_150 <= 16'd881;
      end

      16'd860:
      begin
        register_9 <= register_150;
        program_counter <= 16'd2;
        register_7 <= 16'd861;
      end

      16'd861:
      begin
        register_172 <= register_8;
        register_151 <= 16'd883;
      end

      16'd862:
      begin
        register_9 <= register_151;
        program_counter <= 16'd2;
        register_7 <= 16'd863;
      end

      16'd863:
      begin
        register_172 <= register_8;
        register_16 <= register_112;
        program_counter <= 16'd30;
        register_14 <= 16'd864;
      end

      16'd864:
      begin
        register_172 <= register_15;
        register_152 <= 16'd892;
      end

      16'd865:
      begin
        register_9 <= register_152;
        program_counter <= 16'd2;
        register_7 <= 16'd866;
      end

      16'd866:
      begin
        register_172 <= register_8;
        register_153 <= 16'd894;
      end

      16'd867:
      begin
        register_9 <= register_153;
        program_counter <= 16'd2;
        register_7 <= 16'd868;
      end

      16'd868:
      begin
        register_172 <= register_8;
        register_16 <= register_113;
        program_counter <= 16'd30;
        register_14 <= 16'd869;
      end

      16'd869:
      begin
        register_172 <= register_15;
        register_154 <= 16'd903;
      end

      16'd870:
      begin
        register_9 <= register_154;
        program_counter <= 16'd2;
        register_7 <= 16'd871;
      end

      16'd871:
      begin
        register_172 <= register_8;
        register_155 <= 16'd905;
      end

      16'd872:
      begin
        register_172 <= register_135;
        register_9 <= register_155;
      end

      16'd873:
      begin
        register_172 <= $signed(register_172) + $signed(16'd6);
      end

      16'd874:
      begin
        register_172 <= $signed(register_172) + $signed(register_131);
      end

      16'd875:
      begin
        address <= register_172;
      end

      16'd876:
      begin
        register_172 <= data_out;
      end

      16'd877:
      begin
        register_172 <= data_out;
      end

      16'd878:
      begin
        register_172 <= $signed(register_172) & $signed(16'd1);
      end

      16'd879:
      begin
        register_114 <= register_172;
        register_172 <= register_135;
      end

      16'd880:
      begin
        register_172 <= $signed(register_172) + $signed(16'd6);
      end

      16'd881:
      begin
        register_172 <= $signed(register_172) + $signed(register_131);
      end

      16'd882:
      begin
        address <= register_172;
      end

      16'd883:
      begin
        register_172 <= data_out;
      end

      16'd884:
      begin
        register_172 <= data_out;
      end

      16'd885:
      begin
        register_172 <= $signed(register_172) & $signed(16'd2);
      end

      16'd886:
      begin
        register_115 <= register_172;
        register_172 <= register_135;
      end

      16'd887:
      begin
        register_172 <= $signed(register_172) + $signed(16'd6);
      end

      16'd888:
      begin
        register_172 <= $signed(register_172) + $signed(register_131);
      end

      16'd889:
      begin
        address <= register_172;
      end

      16'd890:
      begin
        register_172 <= data_out;
      end

      16'd891:
      begin
        register_172 <= data_out;
      end

      16'd892:
      begin
        register_172 <= $signed(register_172) & $signed(16'd4);
      end

      16'd893:
      begin
        register_116 <= register_172;
        register_172 <= register_135;
      end

      16'd894:
      begin
        register_172 <= $signed(register_172) + $signed(16'd6);
      end

      16'd895:
      begin
        register_172 <= $signed(register_172) + $signed(register_131);
      end

      16'd896:
      begin
        address <= register_172;
      end

      16'd897:
      begin
        register_172 <= data_out;
      end

      16'd898:
      begin
        register_172 <= data_out;
      end

      16'd899:
      begin
        register_172 <= $signed(register_172) & $signed(16'd8);
      end

      16'd900:
      begin
        register_117 <= register_172;
        register_172 <= register_135;
      end

      16'd901:
      begin
        register_172 <= $signed(register_172) + $signed(16'd6);
      end

      16'd902:
      begin
        register_172 <= $signed(register_172) + $signed(register_131);
      end

      16'd903:
      begin
        address <= register_172;
      end

      16'd904:
      begin
        register_172 <= data_out;
      end

      16'd905:
      begin
        register_172 <= data_out;
      end

      16'd906:
      begin
        register_172 <= $signed(register_172) & $signed(16'd16);
      end

      16'd907:
      begin
        register_118 <= register_172;
        register_172 <= register_135;
      end

      16'd908:
      begin
        register_172 <= $signed(register_172) + $signed(16'd6);
      end

      16'd909:
      begin
        register_172 <= $signed(register_172) + $signed(register_131);
      end

      16'd910:
      begin
        address <= register_172;
      end

      16'd911:
      begin
        register_172 <= data_out;
      end

      16'd912:
      begin
        register_172 <= data_out;
      end

      16'd913:
      begin
        register_172 <= $signed(register_172) & $signed(16'd32);
      end

      16'd914:
      begin
        register_119 <= register_172;
        program_counter <= 16'd2;
        register_7 <= 16'd915;
      end

      16'd915:
      begin
        register_172 <= register_8;
        register_16 <= register_135;
      end

      16'd916:
      begin
        register_16 <= $signed(register_16) + $signed(16'd6);
      end

      16'd917:
      begin
        register_16 <= $signed(register_16) + $signed(register_131);
      end

      16'd918:
      begin
        address <= register_16;
      end

      16'd919:
      begin
        register_16 <= data_out;
      end

      16'd920:
      begin
        register_16 <= data_out;
        program_counter <= 16'd30;
        register_14 <= 16'd921;
      end

      16'd921:
      begin
        register_172 <= register_15;
        register_156 <= 16'd913;
      end

      16'd922:
      begin
        register_9 <= register_156;
        program_counter <= 16'd2;
        register_7 <= 16'd923;
      end

      16'd923:
      begin
        register_172 <= register_8;
        register_130 <= 16'd0;
        program_counter <= register_129;
      end

      16'd924:
      begin
        register_159 <= 16'd915;
        register_160 <= 16'd1939;
        register_161 <= 16'd27;
        register_162 <= 16'd1;
        register_163 <= 16'd2;
        register_164 <= 16'd3;
        register_166 <= 16'd2963;
      end

      16'd925:
      begin
        register_165 <= register_162;
        register_9 <= register_166;
        program_counter <= 16'd2;
        register_7 <= 16'd926;
      end

      16'd926:
      begin
        register_172 <= register_8;
      end

      16'd927:
      begin
        register_172 <= register_165;
        register_173 <= register_162;
      end

      16'd928:
      begin
        register_172 <= $signed(register_172) == $signed(register_173);
      end

      16'd929:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 972;
      end

      16'd930:
      begin
        register_167 <= 16'd2982;
      end

      16'd931:
      begin
        register_9 <= register_167;
        program_counter <= 16'd2;
        register_7 <= 16'd932;
      end

      16'd932:
      begin
        register_172 <= register_8;
        register_131 <= register_159;
        program_counter <= 16'd755;
        register_129 <= 16'd933;
      end

      16'd933:
      begin
        register_172 <= register_130;
      end

      16'd934:
      begin
        register_172 <= register_115;
      end

      16'd935:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 971;
      end

      16'd936:
      begin
        register_168 <= 16'd3006;
      end

      16'd937:
      begin
        register_9 <= register_168;
        program_counter <= 16'd2;
        register_7 <= 16'd938;
      end

      16'd938:
      begin
        register_172 <= register_8;
        register_16 <= 16'd13;
      end

      16'd939:
      begin
        register_16 <= $signed(register_16) + $signed(register_159);
      end

      16'd940:
      begin
        address <= register_16;
      end

      16'd941:
      begin
        register_16 <= data_out;
      end

      16'd942:
      begin
        register_16 <= data_out;
        program_counter <= 16'd30;
        register_14 <= 16'd943;
      end

      16'd943:
      begin
        register_172 <= register_15;
        register_16 <= 16'd14;
      end

      16'd944:
      begin
        register_16 <= $signed(register_16) + $signed(register_159);
      end

      16'd945:
      begin
        address <= register_16;
      end

      16'd946:
      begin
        register_16 <= data_out;
      end

      16'd947:
      begin
        register_16 <= data_out;
        program_counter <= 16'd30;
        register_14 <= 16'd948;
      end

      16'd948:
      begin
        register_172 <= register_15;
        register_169 <= 16'd3034;
      end

      16'd949:
      begin
        register_9 <= register_169;
        program_counter <= 16'd2;
        register_7 <= 16'd950;
      end

      16'd950:
      begin
        register_172 <= register_8;
        register_122 <= register_160;
        register_123 <= 16'd0;
      end

      16'd951:
      begin
        register_172 <= 16'd13;
      end

      16'd952:
      begin
        register_172 <= $signed(register_172) + $signed(register_159);
      end

      16'd953:
      begin
        address <= register_172;
      end

      16'd954:
      begin
        register_172 <= data_out;
      end

      16'd955:
      begin
        register_172 <= data_out;
      end

      16'd956:
      begin
        register_92 <= register_172;
        register_172 <= 16'd14;
      end

      16'd957:
      begin
        register_172 <= $signed(register_172) + $signed(register_159);
      end

      16'd958:
      begin
        address <= register_172;
      end

      16'd959:
      begin
        register_172 <= data_out;
      end

      16'd960:
      begin
        register_172 <= data_out;
      end

      16'd961:
      begin
        register_93 <= register_172;
        register_172 <= register_107;
      end

      16'd962:
      begin
        register_95 <= register_172;
        register_172 <= register_5;
      end

      16'd963:
      begin
        register_94 <= register_172;
        register_172 <= register_110;
      end

      16'd964:
      begin
        register_172 <= $signed(register_172) + $signed(16'd1);
      end

      16'd965:
      begin
        register_99 <= register_172;
        register_172 <= register_109;
      end

      16'd966:
      begin
        register_98 <= register_172;
        register_172 <= 16'd1;
      end

      16'd967:
      begin
        register_102 <= register_172;
        register_172 <= 16'd1;
      end

      16'd968:
      begin
        register_105 <= register_172;
        register_172 <= register_163;
      end

      16'd969:
      begin
        register_165 <= register_172;
        program_counter <= 16'd613;
        register_120 <= 16'd970;
      end

      16'd970:
      begin
        register_172 <= register_121;
        program_counter <= 16'd971;
      end

      16'd971:
      begin
        program_counter <= 16'd991;
      end

      16'd972:
      begin
        register_172 <= register_165;
        register_173 <= register_163;
      end

      16'd973:
      begin
        register_172 <= $signed(register_172) == $signed(register_173);
      end

      16'd974:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 985;
      end

      16'd975:
      begin
        register_170 <= 16'd3036;
      end

      16'd976:
      begin
        register_9 <= register_170;
        program_counter <= 16'd2;
        register_7 <= 16'd977;
      end

      16'd977:
      begin
        register_172 <= register_8;
        register_131 <= register_159;
        program_counter <= 16'd755;
        register_129 <= 16'd978;
      end

      16'd978:
      begin
        register_172 <= register_130;
      end

      16'd979:
      begin
        register_172 <= register_118;
      end

      16'd980:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 984;
      end

      16'd981:
      begin
        register_172 <= register_164;
      end

      16'd982:
      begin
        register_165 <= register_172;
        register_172 <= 16'd0;
      end

      16'd983:
      begin
        register_102 <= register_172;
        program_counter <= 16'd984;
      end

      16'd984:
      begin
        program_counter <= 16'd991;
      end

      16'd985:
      begin
        register_172 <= register_165;
        register_173 <= register_164;
      end

      16'd986:
      begin
        register_172 <= $signed(register_172) == $signed(register_173);
      end

      16'd987:
      begin
        if (register_172 == 16'h0000)
          program_counter <= 991;
      end

      16'd988:
      begin
        register_171 <= 16'd3065;
      end

      16'd989:
      begin
        register_9 <= register_171;
        program_counter <= 16'd2;
        register_7 <= 16'd990;
      end

      16'd990:
      begin
        register_172 <= register_8;
        program_counter <= 16'd991;
      end

      16'd991:
      begin
        program_counter <= 16'd927;
      end

      16'd992:
      begin
        register_172 <= 16'd5;
      end

      16'd993:
      begin
        s_output_leds <= register_172;
        program_counter <= 993;
        s_output_leds_stb <= 1'b1;
        if (s_output_leds_stb == 1'b1 && output_leds_ack == 1'b1) begin
          s_output_leds_stb <= 1'b0;
          program_counter <= 994;
        end
      end

      16'd994:
      begin
        register_172 <= 16'd5;
      end

      16'd995:
      begin
        s_output_checksum <= register_172;
        program_counter <= 995;
        s_output_checksum_stb <= 1'b1;
        if (s_output_checksum_stb == 1'b1 && output_checksum_ack == 1'b1) begin
          s_output_checksum_stb <= 1'b0;
          program_counter <= 996;
        end
      end

      16'd996:
      begin
        register_172 <= input_rs232_rx;
        program_counter <= 996;
        s_input_rs232_rx_ack <= 1'b1;
       if (s_input_rs232_rx_ack == 1'b1 && input_rs232_rx_stb == 1'b1) begin
          s_input_rs232_rx_ack <= 1'b0;
          program_counter <= 16'd997;
        end
      end

      16'd997:
      begin
        register_172 <= input_checksum;
        program_counter <= 997;
        s_input_checksum_ack <= 1'b1;
       if (s_input_checksum_ack == 1'b1 && input_checksum_stb == 1'b1) begin
          s_input_checksum_ack <= 1'b0;
          program_counter <= 16'd998;
        end
      end

      16'd998:
      begin
        register_158 <= 16'd0;
        program_counter <= register_157;
      end

    endcase
    if (rst == 1'b1) begin
      program_counter <= 0;
    end
  end
  assign input_checksum_ack = s_input_checksum_ack;
  assign input_eth_rx_ack = s_input_eth_rx_ack;
  assign input_rs232_rx_ack = s_input_rs232_rx_ack;
  assign output_rs232_tx_stb = s_output_rs232_tx_stb;
  assign output_rs232_tx = s_output_rs232_tx;
  assign output_leds_stb = s_output_leds_stb;
  assign output_leds = s_output_leds;
  assign output_eth_tx_stb = s_output_eth_tx_stb;
  assign output_eth_tx = s_output_eth_tx;
  assign output_checksum_stb = s_output_checksum_stb;
  assign output_checksum = s_output_checksum;

endmodule
