//name : user_design
//tag : c components
//input : input_checksum:16
//input : input_eth_rx:16
//input : input_rs232_rx:16
//output : output_checksum:16
//output : output_leds:16
//output : output_eth_tx:16
//output : output_rs232_tx:16
//source_file : ../source/user_design.c
///User_Design
///===========
///
///*Created by C2CHIP*

  
`timescale 1ns/1ps
module user_design(input_checksum,input_eth_rx,input_rs232_rx,input_checksum_stb,input_eth_rx_stb,input_rs232_rx_stb,output_checksum_ack,output_leds_ack,output_eth_tx_ack,output_rs232_tx_ack,clk,rst,output_checksum,output_leds,output_eth_tx,output_rs232_tx,output_checksum_stb,output_leds_stb,output_eth_tx_stb,output_rs232_tx_stb,input_checksum_ack,input_eth_rx_ack,input_rs232_rx_ack);
  input     [15:0] input_checksum;
  input     [15:0] input_eth_rx;
  input     [15:0] input_rs232_rx;
  input     input_checksum_stb;
  input     input_eth_rx_stb;
  input     input_rs232_rx_stb;
  input     output_checksum_ack;
  input     output_leds_ack;
  input     output_eth_tx_ack;
  input     output_rs232_tx_ack;
  input     clk;
  input     rst;
  output    [15:0] output_checksum;
  output    [15:0] output_leds;
  output    [15:0] output_eth_tx;
  output    [15:0] output_rs232_tx;
  output    output_checksum_stb;
  output    output_leds_stb;
  output    output_eth_tx_stb;
  output    output_rs232_tx_stb;
  output    input_checksum_ack;
  output    input_eth_rx_ack;
  output    input_rs232_rx_ack;
  reg       [15:0] timer;
  reg       [10:0] program_counter;
  reg       [15:0] address;
  reg       [15:0] data_out;
  reg       [15:0] data_in;
  reg       write_enable;
  reg       [15:0] register_0;
  reg       [15:0] register_1;
  reg       [15:0] register_2;
  reg       [15:0] register_3;
  reg       [15:0] register_4;
  reg       [15:0] register_5;
  reg       [15:0] register_6;
  reg       [15:0] register_7;
  reg       [15:0] register_8;
  reg       [15:0] register_9;
  reg       [15:0] register_10;
  reg       [15:0] register_11;
  reg       [15:0] register_12;
  reg       [15:0] register_13;
  reg       [15:0] register_14;
  reg       [15:0] register_15;
  reg       [15:0] register_16;
  reg       [15:0] register_17;
  reg       [15:0] register_18;
  reg       [15:0] register_19;
  reg       [15:0] register_20;
  reg       [15:0] register_21;
  reg       [15:0] register_22;
  reg       [15:0] register_23;
  reg       [15:0] register_24;
  reg       [15:0] register_25;
  reg       [15:0] register_26;
  reg       [15:0] register_27;
  reg       [15:0] register_28;
  reg       [15:0] register_29;
  reg       [15:0] register_30;
  reg       [15:0] register_31;
  reg       [15:0] register_32;
  reg       [15:0] register_33;
  reg       [15:0] register_34;
  reg       [15:0] register_35;
  reg       [15:0] register_36;
  reg       [15:0] register_37;
  reg       [15:0] register_38;
  reg       [15:0] register_39;
  reg       [15:0] register_40;
  reg       [15:0] register_41;
  reg       [15:0] register_42;
  reg       [15:0] register_43;
  reg       [15:0] register_44;
  reg       [15:0] register_45;
  reg       [15:0] register_46;
  reg       [15:0] register_47;
  reg       [15:0] register_48;
  reg       [15:0] register_49;
  reg       [15:0] register_50;
  reg       [15:0] register_51;
  reg       [15:0] register_52;
  reg       [15:0] register_53;
  reg       [15:0] register_54;
  reg       [15:0] register_55;
  reg       [15:0] register_56;
  reg       [15:0] register_57;
  reg       [15:0] register_58;
  reg       [15:0] register_59;
  reg       [15:0] register_60;
  reg       [15:0] register_61;
  reg       [15:0] register_62;
  reg       [15:0] register_63;
  reg       [15:0] register_64;
  reg       [15:0] register_65;
  reg       [15:0] register_66;
  reg       [15:0] register_67;
  reg       [15:0] register_68;
  reg       [15:0] register_69;
  reg       [15:0] register_70;
  reg       [15:0] register_71;
  reg       [15:0] register_72;
  reg       [15:0] register_73;
  reg       [15:0] register_74;
  reg       [15:0] register_75;
  reg       [15:0] register_76;
  reg       [15:0] register_77;
  reg       [15:0] register_78;
  reg       [15:0] register_79;
  reg       [15:0] register_80;
  reg       [15:0] register_81;
  reg       [15:0] register_82;
  reg       [15:0] register_83;
  reg       [15:0] register_84;
  reg       [15:0] register_85;
  reg       [15:0] register_86;
  reg       [15:0] register_87;
  reg       [15:0] register_88;
  reg       [15:0] register_89;
  reg       [15:0] register_90;
  reg       [15:0] register_91;
  reg       [15:0] register_92;
  reg       [15:0] register_93;
  reg       [15:0] register_94;
  reg       [15:0] register_95;
  reg       [15:0] register_96;
  reg       [15:0] register_97;
  reg       [15:0] register_98;
  reg       [15:0] register_99;
  reg       [15:0] register_100;
  reg       [15:0] register_101;
  reg       [15:0] register_102;
  reg       [15:0] register_103;
  reg       [15:0] register_104;
  reg       [15:0] register_105;
  reg       [15:0] register_106;
  reg       [15:0] register_107;
  reg       [15:0] register_108;
  reg       [15:0] register_109;
  reg       [15:0] register_110;
  reg       [15:0] register_111;
  reg       [15:0] register_112;
  reg       [15:0] register_113;
  reg       [15:0] register_114;
  reg       [15:0] register_115;
  reg       [15:0] register_116;
  reg       [15:0] register_117;
  reg       [15:0] register_118;
  reg       [15:0] register_119;
  reg       [15:0] register_120;
  reg       [15:0] register_121;
  reg       [15:0] register_122;
  reg       [15:0] register_123;
  reg       [15:0] register_124;
  reg       [15:0] register_125;
  reg       [15:0] register_126;
  reg       [15:0] register_127;
  reg       [15:0] register_128;
  reg       [15:0] register_129;
  reg       [15:0] register_130;
  reg       [15:0] register_131;
  reg       [15:0] register_132;
  reg       [15:0] register_133;
  reg       [15:0] register_134;
  reg       [15:0] register_135;
  reg       [15:0] register_136;
  reg       [15:0] register_137;
  reg       [15:0] register_138;
  reg       [15:0] register_139;
  reg       [15:0] register_140;
  reg       [15:0] register_141;
  reg       [15:0] register_142;
  reg       [15:0] register_143;
  reg       [15:0] register_144;
  reg       [15:0] register_145;
  reg       [15:0] register_146;
  reg       [15:0] register_147;
  reg       [15:0] register_148;
  reg       [15:0] register_149;
  reg       [15:0] register_150;
  reg       [15:0] register_151;
  reg       [15:0] s_output_checksum_stb;
  reg       [15:0] s_output_leds_stb;
  reg       [15:0] s_output_eth_tx_stb;
  reg       [15:0] s_output_rs232_tx_stb;
  reg       [15:0] s_output_checksum;
  reg       [15:0] s_output_leds;
  reg       [15:0] s_output_eth_tx;
  reg       [15:0] s_output_rs232_tx;
  reg       [15:0] s_input_checksum_ack;
  reg       [15:0] s_input_eth_rx_ack;
  reg       [15:0] s_input_rs232_rx_ack;
  reg [15:0] memory [2693:0];

  //////////////////////////////////////////////////////////////////////////////
  // MEMORY INITIALIZATION                                                      
  //                                                                            
  // In order to reduce program size, array contents have been stored into      
  // memory at initialization. In an FPGA, this will result in the memory being 
  // initialized when the FPGA configures.                                      
  // Memory will not be re-initialized at reset.                                
  // Dissable this behaviour using the no_initialize_memory switch              
  
  initial
  begin
    memory[16'd640] = 16'd111;
    memory[16'd641] = 16'd114;
    memory[16'd642] = 16'd108;
    memory[16'd643] = 16'd100;
    memory[16'd644] = 16'd10;
    memory[16'd645] = 16'd0;
    memory[16'd620] = 16'd77;
    memory[16'd621] = 16'd101;
    memory[16'd622] = 16'd115;
    memory[16'd623] = 16'd115;
    memory[16'd624] = 16'd97;
    memory[16'd625] = 16'd103;
    memory[16'd626] = 16'd101;
    memory[16'd627] = 16'd32;
    memory[16'd628] = 16'd116;
    memory[16'd629] = 16'd111;
    memory[16'd630] = 16'd32;
    memory[16'd631] = 16'd111;
    memory[16'd632] = 16'd117;
    memory[16'd633] = 16'd116;
    memory[16'd634] = 16'd115;
    memory[16'd635] = 16'd105;
    memory[16'd636] = 16'd100;
    memory[16'd637] = 16'd101;
    memory[16'd638] = 16'd32;
    memory[16'd639] = 16'd119;
  end


  //////////////////////////////////////////////////////////////////////////////
  // FSM IMPLEMENTAION OF C PROCESS                                             
  //                                                                            
  // This section of the file contains a Finite State Machine (FSM) implementing
  // the C process. In general execution is sequential, but the compiler will   
  // attempt to execute instructions in parallel if the instruction dependencies
  // allow. Further concurrency can be achieved by executing multiple C         
  // processes concurrently within the device.                                  
  
  always @(posedge clk)
  begin

    if (write_enable == 1'b1) begin
      memory[address] <= data_in;
    end

    data_out <= memory[address];
    write_enable <= 1'b0;
    program_counter <= program_counter + 1;
    timer <= 16'h0000;

    case(program_counter)

      16'd0:
      begin
        register_0 <= 16'd1;
        register_1 <= 16'd515;
        register_2 <= 16'd1029;
        register_3 <= 16'd49320;
        register_4 <= 16'd257;
        register_5 <= 16'd23;
        register_6 <= 16'd0;
        register_7 <= 16'd512;
        register_40 <= 16'd514;
        register_41 <= 16'd530;
        register_42 <= 16'd546;
        register_43 <= 16'd562;
        register_44 <= 16'd578;
        register_45 <= 16'd0;
        register_76 <= 16'd0;
        register_77 <= 16'd0;
        register_78 <= 16'd0;
        register_79 <= 16'd0;
        register_80 <= 16'd610;
        register_81 <= 16'd612;
        register_82 <= 16'd614;
        register_83 <= 16'd1460;
        register_84 <= 16'd0;
        register_85 <= 16'd0;
        register_86 <= 16'd0;
        register_87 <= 16'd0;
        register_88 <= 16'd0;
        register_89 <= 16'd0;
        register_90 <= 16'd0;
        register_91 <= 16'd0;
        register_92 <= 16'd616;
        register_93 <= 16'd618;
        register_94 <= 16'd0;
        register_95 <= 16'd0;
        register_96 <= 16'd0;
        register_97 <= 16'd0;
        register_98 <= 16'd0;
        register_99 <= 16'd0;
        register_100 <= 16'd0;
        register_108 <= 16'd0;
        register_109 <= 16'd0;
        program_counter <= 16'd906;
        register_136 <= 16'd1;
      end

      16'd1:
      begin
        program_counter <= program_counter;
      end

      16'd2:
      begin
        register_150 <= 16'd0;
        register_151 <= 16'd0;
        register_9 <= 16'd0;
      end

      16'd3:
      begin
        register_151 <= $signed(register_151) + $signed(register_7);
      end

      16'd4:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd0;
        register_151 <= 16'd1;
      end

      16'd5:
      begin
        register_151 <= $signed(register_151) + $signed(register_7);
      end

      16'd6:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        program_counter <= register_8;
      end

      16'd7:
      begin
        register_13 <= 16'd0;
        register_150 <= 16'd0;
        register_151 <= register_12;
      end

      16'd8:
      begin
        register_150 <= $signed(register_150) + $signed(register_7);
      end

      16'd9:
      begin
        address <= register_150;
      end

      16'd10:
      begin
        register_150 <= data_out;
      end

      16'd11:
      begin
        register_150 <= data_out;
      end

      16'd12:
      begin
        register_150 <= $signed(register_150) + $signed(register_151);
        register_151 <= register_12;
      end

      16'd13:
      begin
        register_13 <= register_150;
        register_150 <= 16'd0;
      end

      16'd14:
      begin
        register_150 <= $signed(register_150) + $signed(register_7);
      end

      16'd15:
      begin
        address <= register_150;
      end

      16'd16:
      begin
        register_150 <= data_out;
      end

      16'd17:
      begin
        register_150 <= data_out;
      end

      16'd18:
      begin
        register_150 <= $signed(register_150) | $signed(register_151);
      end

      16'd19:
      begin
        register_150 <= $signed(register_150) & $signed(16'd32768);
      end

      16'd20:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 33;
      end

      16'd21:
      begin
        register_150 <= register_13;
      end

      16'd22:
      begin
        register_150 <= $signed(register_150) & $signed(16'd32768);
      end

      16'd23:
      begin
        register_150 <= $signed(register_150) == $signed(16'd0);
      end

      16'd24:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 32;
      end

      16'd25:
      begin
        register_150 <= 16'd1;
        register_151 <= 16'd1;
      end

      16'd26:
      begin
        register_150 <= $signed(register_150) + $signed(register_7);
        register_151 <= $signed(register_151) + $signed(register_7);
      end

      16'd27:
      begin
        address <= register_150;
      end

      16'd28:
      begin
        register_150 <= data_out;
      end

      16'd29:
      begin
        register_150 <= data_out;
      end

      16'd30:
      begin
        register_150 <= $signed(register_150) + $signed(16'd1);
      end

      16'd31:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        program_counter <= 16'd32;
      end

      16'd32:
      begin
        program_counter <= 16'd33;
      end

      16'd33:
      begin
        register_150 <= register_13;
        register_151 <= 16'd0;
        register_11 <= 16'd0;
      end

      16'd34:
      begin
        register_151 <= $signed(register_151) + $signed(register_7);
      end

      16'd35:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        program_counter <= register_10;
      end

      16'd36:
      begin
        register_15 <= 16'd0;
        register_150 <= 16'd1;
      end

      16'd37:
      begin
        register_15 <= $signed(register_15) + $signed(register_7);
        register_150 <= $signed(register_150) + $signed(register_7);
      end

      16'd38:
      begin
        address <= register_15;
      end

      16'd39:
      begin
        register_15 <= data_out;
      end

      16'd40:
      begin
        register_15 <= data_out;
      end

      16'd41:
      begin
        address <= register_150;
      end

      16'd42:
      begin
        register_150 <= data_out;
      end

      16'd43:
      begin
        register_150 <= data_out;
      end

      16'd44:
      begin
        register_15 <= $signed(register_15) + $signed(register_150);
      end

      16'd45:
      begin
        register_15 <= ~register_15;
        program_counter <= register_14;
      end

      16'd46:
      begin
        register_21 <= 16'd0;
        register_22 <= 16'd0;
        register_23 <= 16'd0;
        register_150 <= 16'd0;
        register_151 <= register_20;
      end

      16'd47:
      begin
        register_150 <= $signed(register_150) + $signed(register_19);
      end

      16'd48:
      begin
        address <= register_150;
      end

      16'd49:
      begin
        register_150 <= data_out;
      end

      16'd50:
      begin
        register_150 <= data_out;
      end

      16'd51:
      begin
        register_150 <= $signed(register_150) + $signed(register_151);
        register_151 <= register_20;
      end

      16'd52:
      begin
        register_21 <= register_150;
        register_150 <= 16'd1;
      end

      16'd53:
      begin
        register_150 <= $signed(register_150) + $signed(register_19);
      end

      16'd54:
      begin
        address <= register_150;
      end

      16'd55:
      begin
        register_150 <= data_out;
      end

      16'd56:
      begin
        register_150 <= data_out;
      end

      16'd57:
      begin
        register_22 <= register_150;
        register_150 <= 16'd0;
      end

      16'd58:
      begin
        register_150 <= $signed(register_150) + $signed(register_19);
      end

      16'd59:
      begin
        address <= register_150;
      end

      16'd60:
      begin
        register_150 <= data_out;
      end

      16'd61:
      begin
        register_150 <= data_out;
      end

      16'd62:
      begin
        register_150 <= $signed(register_150) | $signed(register_151);
      end

      16'd63:
      begin
        register_150 <= $signed(register_150) & $signed(16'd32768);
      end

      16'd64:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 73;
      end

      16'd65:
      begin
        register_150 <= register_21;
      end

      16'd66:
      begin
        register_150 <= $signed(register_150) & $signed(16'd32768);
      end

      16'd67:
      begin
        register_150 <= $signed(register_150) == $signed(16'd0);
      end

      16'd68:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 72;
      end

      16'd69:
      begin
        register_150 <= register_22;
      end

      16'd70:
      begin
        register_150 <= $signed(register_150) + $signed(16'd1);
      end

      16'd71:
      begin
        register_22 <= register_150;
        program_counter <= 16'd72;
      end

      16'd72:
      begin
        program_counter <= 16'd73;
      end

      16'd73:
      begin
        register_150 <= register_21;
        register_151 <= 16'd0;
      end

      16'd74:
      begin
        register_151 <= $signed(register_151) + $signed(register_18);
      end

      16'd75:
      begin
        address <= register_151;
      end

      16'd76:
      begin
        register_151 <= data_out;
      end

      16'd77:
      begin
        register_151 <= data_out;
      end

      16'd78:
      begin
        register_150 <= $signed(register_150) != $signed(register_151);
      end

      16'd79:
      begin
        if (register_150 != 16'h0000)
          program_counter <= 16'd86;
      end

      16'd80:
      begin
        register_150 <= register_22;
        register_151 <= 16'd1;
      end

      16'd81:
      begin
        register_151 <= $signed(register_151) + $signed(register_18);
      end

      16'd82:
      begin
        address <= register_151;
      end

      16'd83:
      begin
        register_151 <= data_out;
      end

      16'd84:
      begin
        register_151 <= data_out;
      end

      16'd85:
      begin
        register_150 <= $signed(register_150) != $signed(register_151);
      end

      16'd86:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 93;
      end

      16'd87:
      begin
        register_150 <= register_21;
        register_151 <= 16'd0;
      end

      16'd88:
      begin
        register_151 <= $signed(register_151) + $signed(register_18);
      end

      16'd89:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_22;
        register_151 <= 16'd1;
      end

      16'd90:
      begin
        register_151 <= $signed(register_151) + $signed(register_18);
      end

      16'd91:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd1;
      end

      16'd92:
      begin
        register_23 <= register_150;
        program_counter <= 16'd93;
      end

      16'd93:
      begin
        register_17 <= register_23;
        program_counter <= register_16;
      end

      16'd94:
      begin
        register_32 <= 16'd0;
        register_33 <= 16'd0;
        register_150 <= register_28;
        register_151 <= 16'd0;
      end

      16'd95:
      begin
        register_151 <= $signed(register_151) + $signed(register_26);
      end

      16'd96:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_29;
        register_151 <= 16'd1;
      end

      16'd97:
      begin
        register_151 <= $signed(register_151) + $signed(register_26);
      end

      16'd98:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_30;
        register_151 <= 16'd2;
      end

      16'd99:
      begin
        register_151 <= $signed(register_151) + $signed(register_26);
      end

      16'd100:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_0;
        register_151 <= 16'd3;
      end

      16'd101:
      begin
        register_151 <= $signed(register_151) + $signed(register_26);
      end

      16'd102:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_1;
        register_151 <= 16'd4;
      end

      16'd103:
      begin
        register_151 <= $signed(register_151) + $signed(register_26);
      end

      16'd104:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_2;
        register_151 <= 16'd5;
      end

      16'd105:
      begin
        register_151 <= $signed(register_151) + $signed(register_26);
      end

      16'd106:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_31;
        register_151 <= 16'd6;
      end

      16'd107:
      begin
        register_151 <= $signed(register_151) + $signed(register_26);
      end

      16'd108:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_27;
      end

      16'd109:
      begin
        s_output_eth_tx <= register_150;
        program_counter <= 109;
        s_output_eth_tx_stb <= 1'b1;
        if (s_output_eth_tx_stb == 1'b1 && output_eth_tx_ack == 1'b1) begin
          s_output_eth_tx_stb <= 1'b0;
          program_counter <= 110;
        end
      end

      16'd110:
      begin
        register_150 <= 16'd0;
      end

      16'd111:
      begin
        register_33 <= register_150;
        register_150 <= 16'd0;
      end

      16'd112:
      begin
        register_32 <= register_150;
      end

      16'd113:
      begin
        register_150 <= register_32;
        register_151 <= register_27;
      end

      16'd114:
      begin
        register_150 <= $signed(register_150) < $signed(register_151);
      end

      16'd115:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 128;
      end

      16'd116:
      begin
        register_150 <= register_33;
      end

      16'd117:
      begin
        register_150 <= $signed(register_150) + $signed(register_26);
      end

      16'd118:
      begin
        address <= register_150;
      end

      16'd119:
      begin
        register_150 <= data_out;
      end

      16'd120:
      begin
        register_150 <= data_out;
      end

      16'd121:
      begin
        s_output_eth_tx <= register_150;
        program_counter <= 121;
        s_output_eth_tx_stb <= 1'b1;
        if (s_output_eth_tx_stb == 1'b1 && output_eth_tx_ack == 1'b1) begin
          s_output_eth_tx_stb <= 1'b0;
          program_counter <= 122;
        end
      end

      16'd122:
      begin
        register_150 <= register_33;
      end

      16'd123:
      begin
        register_150 <= $signed(register_150) + $signed(16'd1);
      end

      16'd124:
      begin
        register_33 <= register_150;
      end

      16'd125:
      begin
        register_150 <= register_32;
      end

      16'd126:
      begin
        register_150 <= $signed(register_150) + $signed(16'd2);
      end

      16'd127:
      begin
        register_32 <= register_150;
        program_counter <= 16'd113;
      end

      16'd128:
      begin
        register_25 <= 16'd0;
        program_counter <= register_24;
      end

      16'd129:
      begin
        register_37 <= 16'd0;
        register_38 <= 16'd0;
        register_39 <= 16'd0;
      end

      16'd130:
      begin
        register_150 <= input_eth_rx;
        program_counter <= 130;
        s_input_eth_rx_ack <= 1'b1;
       if (s_input_eth_rx_ack == 1'b1 && input_eth_rx_stb == 1'b1) begin
          s_input_eth_rx_ack <= 1'b0;
          program_counter <= 16'd131;
        end
      end

      16'd131:
      begin
        register_37 <= register_150;
        register_150 <= 16'd0;
      end

      16'd132:
      begin
        register_38 <= register_150;
        register_150 <= 16'd0;
      end

      16'd133:
      begin
        register_39 <= register_150;
      end

      16'd134:
      begin
        register_150 <= register_39;
        register_151 <= register_37;
      end

      16'd135:
      begin
        register_150 <= $signed(register_150) < $signed(register_151);
      end

      16'd136:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 146;
      end

      16'd137:
      begin
        register_150 <= input_eth_rx;
        program_counter <= 137;
        s_input_eth_rx_ack <= 1'b1;
       if (s_input_eth_rx_ack == 1'b1 && input_eth_rx_stb == 1'b1) begin
          s_input_eth_rx_ack <= 1'b0;
          program_counter <= 16'd138;
        end
      end

      16'd138:
      begin
        register_151 <= register_38;
      end

      16'd139:
      begin
        register_151 <= $signed(register_151) + $signed(register_36);
      end

      16'd140:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_38;
      end

      16'd141:
      begin
        register_150 <= $signed(register_150) + $signed(16'd1);
      end

      16'd142:
      begin
        register_38 <= register_150;
      end

      16'd143:
      begin
        register_150 <= register_39;
      end

      16'd144:
      begin
        register_150 <= $signed(register_150) + $signed(16'd2);
      end

      16'd145:
      begin
        register_39 <= register_150;
        program_counter <= 16'd134;
      end

      16'd146:
      begin
        register_150 <= 16'd0;
        register_151 <= register_0;
      end

      16'd147:
      begin
        register_150 <= $signed(register_150) + $signed(register_36);
      end

      16'd148:
      begin
        address <= register_150;
      end

      16'd149:
      begin
        register_150 <= data_out;
      end

      16'd150:
      begin
        register_150 <= data_out;
      end

      16'd151:
      begin
        register_150 <= $signed(register_150) != $signed(register_151);
      end

      16'd152:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 159;
      end

      16'd153:
      begin
        register_150 <= 16'd0;
      end

      16'd154:
      begin
        register_150 <= $signed(register_150) + $signed(register_36);
      end

      16'd155:
      begin
        address <= register_150;
      end

      16'd156:
      begin
        register_150 <= data_out;
      end

      16'd157:
      begin
        register_150 <= data_out;
      end

      16'd158:
      begin
        register_150 <= $signed(register_150) != $signed(16'd65535);
      end

      16'd159:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 162;
      end

      16'd160:
      begin
        program_counter <= 16'd130;
      end

      16'd161:
      begin
        program_counter <= 16'd162;
      end

      16'd162:
      begin
        register_150 <= 16'd1;
        register_151 <= register_1;
      end

      16'd163:
      begin
        register_150 <= $signed(register_150) + $signed(register_36);
      end

      16'd164:
      begin
        address <= register_150;
      end

      16'd165:
      begin
        register_150 <= data_out;
      end

      16'd166:
      begin
        register_150 <= data_out;
      end

      16'd167:
      begin
        register_150 <= $signed(register_150) != $signed(register_151);
      end

      16'd168:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 175;
      end

      16'd169:
      begin
        register_150 <= 16'd1;
      end

      16'd170:
      begin
        register_150 <= $signed(register_150) + $signed(register_36);
      end

      16'd171:
      begin
        address <= register_150;
      end

      16'd172:
      begin
        register_150 <= data_out;
      end

      16'd173:
      begin
        register_150 <= data_out;
      end

      16'd174:
      begin
        register_150 <= $signed(register_150) != $signed(16'd65535);
      end

      16'd175:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 178;
      end

      16'd176:
      begin
        program_counter <= 16'd130;
      end

      16'd177:
      begin
        program_counter <= 16'd178;
      end

      16'd178:
      begin
        register_150 <= 16'd2;
        register_151 <= register_2;
      end

      16'd179:
      begin
        register_150 <= $signed(register_150) + $signed(register_36);
      end

      16'd180:
      begin
        address <= register_150;
      end

      16'd181:
      begin
        register_150 <= data_out;
      end

      16'd182:
      begin
        register_150 <= data_out;
      end

      16'd183:
      begin
        register_150 <= $signed(register_150) != $signed(register_151);
      end

      16'd184:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 191;
      end

      16'd185:
      begin
        register_150 <= 16'd2;
      end

      16'd186:
      begin
        register_150 <= $signed(register_150) + $signed(register_36);
      end

      16'd187:
      begin
        address <= register_150;
      end

      16'd188:
      begin
        register_150 <= data_out;
      end

      16'd189:
      begin
        register_150 <= data_out;
      end

      16'd190:
      begin
        register_150 <= $signed(register_150) != $signed(16'd65535);
      end

      16'd191:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 194;
      end

      16'd192:
      begin
        program_counter <= 16'd130;
      end

      16'd193:
      begin
        program_counter <= 16'd194;
      end

      16'd194:
      begin
        register_150 <= 16'd6;
      end

      16'd195:
      begin
        register_150 <= $signed(register_150) + $signed(register_36);
      end

      16'd196:
      begin
        address <= register_150;
      end

      16'd197:
      begin
        register_150 <= data_out;
      end

      16'd198:
      begin
        register_150 <= data_out;
      end

      16'd199:
      begin
        register_150 <= $signed(register_150) == $signed(16'd2054);
      end

      16'd200:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 264;
      end

      16'd201:
      begin
        register_150 <= 16'd10;
      end

      16'd202:
      begin
        register_150 <= $signed(register_150) + $signed(register_36);
      end

      16'd203:
      begin
        address <= register_150;
      end

      16'd204:
      begin
        register_150 <= data_out;
      end

      16'd205:
      begin
        register_150 <= data_out;
      end

      16'd206:
      begin
        register_150 <= $signed(register_150) == $signed(16'd1);
      end

      16'd207:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 262;
      end

      16'd208:
      begin
        register_150 <= 16'd1;
        register_151 <= 16'd7;
        register_26 <= register_6;
        register_27 <= 16'd64;
        register_28 <= 16'd11;
        register_29 <= 16'd12;
        register_30 <= 16'd13;
        register_31 <= 16'd2054;
      end

      16'd209:
      begin
        register_151 <= $signed(register_151) + $signed(register_6);
        register_28 <= $signed(register_28) + $signed(register_36);
        register_29 <= $signed(register_29) + $signed(register_36);
        register_30 <= $signed(register_30) + $signed(register_36);
      end

      16'd210:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd2048;
        register_151 <= 16'd8;
      end

      16'd211:
      begin
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd212:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd1540;
        register_151 <= 16'd9;
      end

      16'd213:
      begin
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd214:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd2;
        register_151 <= 16'd10;
      end

      16'd215:
      begin
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd216:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_0;
        register_151 <= 16'd11;
      end

      16'd217:
      begin
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd218:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_1;
        register_151 <= 16'd12;
      end

      16'd219:
      begin
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd220:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_2;
        register_151 <= 16'd13;
      end

      16'd221:
      begin
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd222:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_3;
        register_151 <= 16'd14;
      end

      16'd223:
      begin
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd224:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_4;
        register_151 <= 16'd15;
      end

      16'd225:
      begin
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd226:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd11;
        register_151 <= 16'd16;
      end

      16'd227:
      begin
        register_150 <= $signed(register_150) + $signed(register_36);
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd228:
      begin
        address <= register_150;
      end

      16'd229:
      begin
        register_150 <= data_out;
      end

      16'd230:
      begin
        register_150 <= data_out;
      end

      16'd231:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd12;
        register_151 <= 16'd17;
      end

      16'd232:
      begin
        register_150 <= $signed(register_150) + $signed(register_36);
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd233:
      begin
        address <= register_150;
      end

      16'd234:
      begin
        register_150 <= data_out;
      end

      16'd235:
      begin
        register_150 <= data_out;
      end

      16'd236:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd13;
        register_151 <= 16'd18;
      end

      16'd237:
      begin
        register_150 <= $signed(register_150) + $signed(register_36);
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd238:
      begin
        address <= register_150;
      end

      16'd239:
      begin
        register_150 <= data_out;
      end

      16'd240:
      begin
        register_150 <= data_out;
      end

      16'd241:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd14;
        register_151 <= 16'd19;
      end

      16'd242:
      begin
        register_150 <= $signed(register_150) + $signed(register_36);
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd243:
      begin
        address <= register_150;
      end

      16'd244:
      begin
        register_150 <= data_out;
      end

      16'd245:
      begin
        register_150 <= data_out;
      end

      16'd246:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd15;
        register_151 <= 16'd20;
      end

      16'd247:
      begin
        register_150 <= $signed(register_150) + $signed(register_36);
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd248:
      begin
        address <= register_150;
      end

      16'd249:
      begin
        register_150 <= data_out;
      end

      16'd250:
      begin
        register_150 <= data_out;
      end

      16'd251:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
      end

      16'd252:
      begin
        address <= register_28;
      end

      16'd253:
      begin
        register_28 <= data_out;
      end

      16'd254:
      begin
        register_28 <= data_out;
      end

      16'd255:
      begin
        address <= register_29;
      end

      16'd256:
      begin
        register_29 <= data_out;
      end

      16'd257:
      begin
        register_29 <= data_out;
      end

      16'd258:
      begin
        address <= register_30;
      end

      16'd259:
      begin
        register_30 <= data_out;
      end

      16'd260:
      begin
        register_30 <= data_out;
        program_counter <= 16'd94;
        register_24 <= 16'd261;
      end

      16'd261:
      begin
        register_150 <= register_25;
        program_counter <= 16'd262;
      end

      16'd262:
      begin
        program_counter <= 16'd130;
      end

      16'd263:
      begin
        program_counter <= 16'd264;
      end

      16'd264:
      begin
        program_counter <= 16'd266;
      end

      16'd265:
      begin
        program_counter <= 16'd130;
      end

      16'd266:
      begin
        register_35 <= register_37;
        program_counter <= register_34;
      end

      16'd267:
      begin
        register_50 <= 16'd0;
        register_51 <= 16'd0;
        register_52 <= 16'd594;
        register_53 <= 16'd0;
        register_150 <= 16'd0;
      end

      16'd268:
      begin
        register_53 <= register_150;
      end

      16'd269:
      begin
        register_150 <= register_53;
      end

      16'd270:
      begin
        register_150 <= $signed(register_150) < $signed(16'd16);
      end

      16'd271:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 291;
      end

      16'd272:
      begin
        register_150 <= register_53;
        register_151 <= register_48;
      end

      16'd273:
      begin
        register_150 <= $signed(register_150) + $signed(register_40);
      end

      16'd274:
      begin
        address <= register_150;
      end

      16'd275:
      begin
        register_150 <= data_out;
      end

      16'd276:
      begin
        register_150 <= data_out;
      end

      16'd277:
      begin
        register_150 <= $signed(register_150) == $signed(register_151);
      end

      16'd278:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 285;
      end

      16'd279:
      begin
        register_150 <= register_53;
        register_151 <= register_49;
      end

      16'd280:
      begin
        register_150 <= $signed(register_150) + $signed(register_41);
      end

      16'd281:
      begin
        address <= register_150;
      end

      16'd282:
      begin
        register_150 <= data_out;
      end

      16'd283:
      begin
        register_150 <= data_out;
      end

      16'd284:
      begin
        register_150 <= $signed(register_150) == $signed(register_151);
      end

      16'd285:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 288;
      end

      16'd286:
      begin
        register_47 <= register_53;
        program_counter <= register_46;
      end

      16'd287:
      begin
        program_counter <= 16'd288;
      end

      16'd288:
      begin
        register_150 <= register_53;
      end

      16'd289:
      begin
        register_150 <= $signed(register_150) + $signed(16'd1);
      end

      16'd290:
      begin
        register_53 <= register_150;
        program_counter <= 16'd269;
      end

      16'd291:
      begin
        register_150 <= 16'd1;
        register_151 <= 16'd7;
        register_26 <= register_6;
        register_27 <= 16'd64;
        register_28 <= 16'd65535;
        register_29 <= 16'd65535;
        register_30 <= 16'd65535;
        register_31 <= 16'd2054;
      end

      16'd292:
      begin
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd293:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd2048;
        register_151 <= 16'd8;
      end

      16'd294:
      begin
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd295:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd1540;
        register_151 <= 16'd9;
      end

      16'd296:
      begin
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd297:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd1;
        register_151 <= 16'd10;
      end

      16'd298:
      begin
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd299:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_0;
        register_151 <= 16'd11;
      end

      16'd300:
      begin
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd301:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_1;
        register_151 <= 16'd12;
      end

      16'd302:
      begin
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd303:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_2;
        register_151 <= 16'd13;
      end

      16'd304:
      begin
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd305:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_3;
        register_151 <= 16'd14;
      end

      16'd306:
      begin
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd307:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_4;
        register_151 <= 16'd15;
      end

      16'd308:
      begin
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd309:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_48;
        register_151 <= 16'd19;
      end

      16'd310:
      begin
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd311:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_49;
        register_151 <= 16'd20;
      end

      16'd312:
      begin
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd313:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        program_counter <= 16'd94;
        register_24 <= 16'd314;
      end

      16'd314:
      begin
        register_150 <= register_25;
      end

      16'd315:
      begin
        register_150 <= input_eth_rx;
        program_counter <= 315;
        s_input_eth_rx_ack <= 1'b1;
       if (s_input_eth_rx_ack == 1'b1 && input_eth_rx_stb == 1'b1) begin
          s_input_eth_rx_ack <= 1'b0;
          program_counter <= 16'd316;
        end
      end

      16'd316:
      begin
        register_50 <= register_150;
        register_150 <= 16'd0;
      end

      16'd317:
      begin
        register_53 <= register_150;
        register_150 <= 16'd0;
      end

      16'd318:
      begin
        register_51 <= register_150;
      end

      16'd319:
      begin
        register_150 <= register_51;
        register_151 <= register_50;
      end

      16'd320:
      begin
        register_150 <= $signed(register_150) < $signed(register_151);
      end

      16'd321:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 336;
      end

      16'd322:
      begin
        register_150 <= register_53;
      end

      16'd323:
      begin
        register_150 <= $signed(register_150) < $signed(16'd16);
      end

      16'd324:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 329;
      end

      16'd325:
      begin
        register_150 <= input_eth_rx;
        program_counter <= 325;
        s_input_eth_rx_ack <= 1'b1;
       if (s_input_eth_rx_ack == 1'b1 && input_eth_rx_stb == 1'b1) begin
          s_input_eth_rx_ack <= 1'b0;
          program_counter <= 16'd326;
        end
      end

      16'd326:
      begin
        register_151 <= register_53;
      end

      16'd327:
      begin
        register_151 <= $signed(register_151) + $signed(register_52);
      end

      16'd328:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        program_counter <= 16'd330;
      end

      16'd329:
      begin
        register_150 <= input_eth_rx;
        program_counter <= 329;
        s_input_eth_rx_ack <= 1'b1;
       if (s_input_eth_rx_ack == 1'b1 && input_eth_rx_stb == 1'b1) begin
          s_input_eth_rx_ack <= 1'b0;
          program_counter <= 16'd330;
        end
      end

      16'd330:
      begin
        register_150 <= register_53;
      end

      16'd331:
      begin
        register_150 <= $signed(register_150) + $signed(16'd1);
      end

      16'd332:
      begin
        register_53 <= register_150;
      end

      16'd333:
      begin
        register_150 <= register_51;
      end

      16'd334:
      begin
        register_150 <= $signed(register_150) + $signed(16'd2);
      end

      16'd335:
      begin
        register_51 <= register_150;
        program_counter <= 16'd319;
      end

      16'd336:
      begin
        register_150 <= 16'd6;
      end

      16'd337:
      begin
        register_150 <= $signed(register_150) + $signed(register_52);
      end

      16'd338:
      begin
        address <= register_150;
      end

      16'd339:
      begin
        register_150 <= data_out;
      end

      16'd340:
      begin
        register_150 <= data_out;
      end

      16'd341:
      begin
        register_150 <= $signed(register_150) == $signed(16'd2054);
      end

      16'd342:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 349;
      end

      16'd343:
      begin
        register_150 <= 16'd10;
      end

      16'd344:
      begin
        register_150 <= $signed(register_150) + $signed(register_52);
      end

      16'd345:
      begin
        address <= register_150;
      end

      16'd346:
      begin
        register_150 <= data_out;
      end

      16'd347:
      begin
        register_150 <= data_out;
      end

      16'd348:
      begin
        register_150 <= $signed(register_150) == $signed(16'd2);
      end

      16'd349:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 395;
      end

      16'd350:
      begin
        register_150 <= 16'd14;
        register_151 <= register_48;
      end

      16'd351:
      begin
        register_150 <= $signed(register_150) + $signed(register_52);
      end

      16'd352:
      begin
        address <= register_150;
      end

      16'd353:
      begin
        register_150 <= data_out;
      end

      16'd354:
      begin
        register_150 <= data_out;
      end

      16'd355:
      begin
        register_150 <= $signed(register_150) == $signed(register_151);
      end

      16'd356:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 363;
      end

      16'd357:
      begin
        register_150 <= 16'd15;
        register_151 <= register_49;
      end

      16'd358:
      begin
        register_150 <= $signed(register_150) + $signed(register_52);
      end

      16'd359:
      begin
        address <= register_150;
      end

      16'd360:
      begin
        register_150 <= data_out;
      end

      16'd361:
      begin
        register_150 <= data_out;
      end

      16'd362:
      begin
        register_150 <= $signed(register_150) == $signed(register_151);
      end

      16'd363:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 394;
      end

      16'd364:
      begin
        register_150 <= register_48;
        register_151 <= register_45;
      end

      16'd365:
      begin
        register_151 <= $signed(register_151) + $signed(register_40);
      end

      16'd366:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_49;
        register_151 <= register_45;
      end

      16'd367:
      begin
        register_151 <= $signed(register_151) + $signed(register_41);
      end

      16'd368:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd11;
        register_151 <= register_45;
      end

      16'd369:
      begin
        register_150 <= $signed(register_150) + $signed(register_52);
        register_151 <= $signed(register_151) + $signed(register_42);
      end

      16'd370:
      begin
        address <= register_150;
      end

      16'd371:
      begin
        register_150 <= data_out;
      end

      16'd372:
      begin
        register_150 <= data_out;
      end

      16'd373:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd12;
        register_151 <= register_45;
      end

      16'd374:
      begin
        register_150 <= $signed(register_150) + $signed(register_52);
        register_151 <= $signed(register_151) + $signed(register_43);
      end

      16'd375:
      begin
        address <= register_150;
      end

      16'd376:
      begin
        register_150 <= data_out;
      end

      16'd377:
      begin
        register_150 <= data_out;
      end

      16'd378:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd13;
        register_151 <= register_45;
      end

      16'd379:
      begin
        register_150 <= $signed(register_150) + $signed(register_52);
        register_151 <= $signed(register_151) + $signed(register_44);
      end

      16'd380:
      begin
        address <= register_150;
      end

      16'd381:
      begin
        register_150 <= data_out;
      end

      16'd382:
      begin
        register_150 <= data_out;
      end

      16'd383:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_45;
      end

      16'd384:
      begin
        register_53 <= register_150;
        register_150 <= register_45;
      end

      16'd385:
      begin
        register_150 <= $signed(register_150) + $signed(16'd1);
      end

      16'd386:
      begin
        register_45 <= register_150;
      end

      16'd387:
      begin
        register_150 <= register_45;
      end

      16'd388:
      begin
        register_150 <= $signed(register_150) == $signed(16'd16);
      end

      16'd389:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 392;
      end

      16'd390:
      begin
        register_150 <= 16'd0;
      end

      16'd391:
      begin
        register_45 <= register_150;
        program_counter <= 16'd392;
      end

      16'd392:
      begin
        register_47 <= register_53;
        program_counter <= register_46;
      end

      16'd393:
      begin
        program_counter <= 16'd394;
      end

      16'd394:
      begin
        program_counter <= 16'd395;
      end

      16'd395:
      begin
        program_counter <= 16'd315;
      end

      16'd396:
      begin
        register_61 <= 16'd0;
        register_62 <= 16'd0;
        register_63 <= 16'd0;
        register_48 <= register_59;
        register_49 <= register_60;
        program_counter <= 16'd267;
        register_46 <= 16'd397;
      end

      16'd397:
      begin
        register_150 <= register_47;
        register_151 <= 16'd7;
      end

      16'd398:
      begin
        register_63 <= register_150;
        register_150 <= 16'd17664;
        register_151 <= $signed(register_151) + $signed(register_56);
      end

      16'd399:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_57;
        register_151 <= 16'd8;
      end

      16'd400:
      begin
        register_151 <= $signed(register_151) + $signed(register_56);
      end

      16'd401:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd0;
        register_151 <= 16'd9;
      end

      16'd402:
      begin
        register_151 <= $signed(register_151) + $signed(register_56);
      end

      16'd403:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd16384;
        register_151 <= 16'd10;
      end

      16'd404:
      begin
        register_151 <= $signed(register_151) + $signed(register_56);
      end

      16'd405:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_58;
        register_151 <= 16'd11;
      end

      16'd406:
      begin
        register_150 <= $signed(16'd65280) | $signed(register_150);
        register_151 <= $signed(register_151) + $signed(register_56);
      end

      16'd407:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd0;
        register_151 <= 16'd12;
      end

      16'd408:
      begin
        register_151 <= $signed(register_151) + $signed(register_56);
      end

      16'd409:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_3;
        register_151 <= 16'd13;
      end

      16'd410:
      begin
        register_151 <= $signed(register_151) + $signed(register_56);
      end

      16'd411:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_4;
        register_151 <= 16'd14;
      end

      16'd412:
      begin
        register_151 <= $signed(register_151) + $signed(register_56);
      end

      16'd413:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_59;
        register_151 <= 16'd15;
      end

      16'd414:
      begin
        register_151 <= $signed(register_151) + $signed(register_56);
      end

      16'd415:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_60;
        register_151 <= 16'd16;
      end

      16'd416:
      begin
        register_151 <= $signed(register_151) + $signed(register_56);
      end

      16'd417:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_57;
      end

      16'd418:
      begin
        register_150 <= $signed(register_150) + $signed(16'd14);
      end

      16'd419:
      begin
        register_61 <= register_150;
        program_counter <= 16'd2;
        register_8 <= 16'd420;
      end

      16'd420:
      begin
        register_150 <= register_9;
      end

      16'd421:
      begin
        register_150 <= 16'd7;
      end

      16'd422:
      begin
        register_62 <= register_150;
      end

      16'd423:
      begin
        register_150 <= register_62;
      end

      16'd424:
      begin
        register_150 <= $signed(register_150) <= $signed(16'd16);
      end

      16'd425:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 435;
      end

      16'd426:
      begin
        register_12 <= register_62;
      end

      16'd427:
      begin
        register_12 <= $signed(register_12) + $signed(register_56);
      end

      16'd428:
      begin
        address <= register_12;
      end

      16'd429:
      begin
        register_12 <= data_out;
      end

      16'd430:
      begin
        register_12 <= data_out;
        program_counter <= 16'd7;
        register_10 <= 16'd431;
      end

      16'd431:
      begin
        register_150 <= register_11;
      end

      16'd432:
      begin
        register_150 <= register_62;
      end

      16'd433:
      begin
        register_150 <= $signed(register_150) + $signed(16'd1);
      end

      16'd434:
      begin
        register_62 <= register_150;
        program_counter <= 16'd423;
      end

      16'd435:
      begin
        program_counter <= 16'd36;
        register_14 <= 16'd436;
      end

      16'd436:
      begin
        register_150 <= register_15;
        register_151 <= 16'd12;
      end

      16'd437:
      begin
        register_151 <= $signed(register_151) + $signed(register_56);
      end

      16'd438:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_61;
      end

      16'd439:
      begin
        register_150 <= $signed(register_150) < $signed(16'd64);
      end

      16'd440:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 443;
      end

      16'd441:
      begin
        register_150 <= 16'd64;
      end

      16'd442:
      begin
        register_61 <= register_150;
        program_counter <= 16'd443;
      end

      16'd443:
      begin
        register_26 <= register_56;
        register_27 <= register_61;
        register_28 <= register_63;
        register_29 <= register_63;
        register_30 <= register_63;
        register_31 <= 16'd2048;
      end

      16'd444:
      begin
        register_28 <= $signed(register_28) + $signed(register_42);
        register_29 <= $signed(register_29) + $signed(register_43);
        register_30 <= $signed(register_30) + $signed(register_44);
      end

      16'd445:
      begin
        address <= register_28;
      end

      16'd446:
      begin
        register_28 <= data_out;
      end

      16'd447:
      begin
        register_28 <= data_out;
      end

      16'd448:
      begin
        address <= register_29;
      end

      16'd449:
      begin
        register_29 <= data_out;
      end

      16'd450:
      begin
        register_29 <= data_out;
      end

      16'd451:
      begin
        address <= register_30;
      end

      16'd452:
      begin
        register_30 <= data_out;
      end

      16'd453:
      begin
        register_30 <= data_out;
        program_counter <= 16'd94;
        register_24 <= 16'd454;
      end

      16'd454:
      begin
        register_150 <= register_25;
        register_55 <= 16'd0;
        program_counter <= register_54;
      end

      16'd455:
      begin
        register_67 <= 16'd0;
        register_68 <= 16'd0;
        register_69 <= 16'd0;
        register_70 <= 16'd0;
        register_71 <= 16'd0;
        register_72 <= 16'd0;
        register_73 <= 16'd0;
        register_74 <= 16'd0;
        register_75 <= 16'd0;
      end

      16'd456:
      begin
        register_36 <= register_66;
        program_counter <= 16'd129;
        register_34 <= 16'd457;
      end

      16'd457:
      begin
        register_150 <= register_35;
      end

      16'd458:
      begin
        register_61 <= register_150;
        register_150 <= 16'd6;
      end

      16'd459:
      begin
        register_150 <= $signed(register_150) + $signed(register_66);
      end

      16'd460:
      begin
        address <= register_150;
      end

      16'd461:
      begin
        register_150 <= data_out;
      end

      16'd462:
      begin
        register_150 <= data_out;
      end

      16'd463:
      begin
        register_150 <= $signed(register_150) == $signed(16'd2048);
      end

      16'd464:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 578;
      end

      16'd465:
      begin
        register_150 <= 16'd15;
        register_151 <= register_3;
      end

      16'd466:
      begin
        register_150 <= $signed(register_150) + $signed(register_66);
      end

      16'd467:
      begin
        address <= register_150;
      end

      16'd468:
      begin
        register_150 <= data_out;
      end

      16'd469:
      begin
        register_150 <= data_out;
      end

      16'd470:
      begin
        register_150 <= $signed(register_150) != $signed(register_151);
      end

      16'd471:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 474;
      end

      16'd472:
      begin
        program_counter <= 16'd456;
      end

      16'd473:
      begin
        program_counter <= 16'd474;
      end

      16'd474:
      begin
        register_150 <= 16'd16;
        register_151 <= register_4;
      end

      16'd475:
      begin
        register_150 <= $signed(register_150) + $signed(register_66);
      end

      16'd476:
      begin
        address <= register_150;
      end

      16'd477:
      begin
        register_150 <= data_out;
      end

      16'd478:
      begin
        register_150 <= data_out;
      end

      16'd479:
      begin
        register_150 <= $signed(register_150) != $signed(register_151);
      end

      16'd480:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 483;
      end

      16'd481:
      begin
        program_counter <= 16'd456;
      end

      16'd482:
      begin
        program_counter <= 16'd483;
      end

      16'd483:
      begin
        register_150 <= 16'd11;
      end

      16'd484:
      begin
        register_150 <= $signed(register_150) + $signed(register_66);
      end

      16'd485:
      begin
        address <= register_150;
      end

      16'd486:
      begin
        register_150 <= data_out;
      end

      16'd487:
      begin
        register_150 <= data_out;
      end

      16'd488:
      begin
        register_150 <= $signed(register_150) & $signed(16'd255);
      end

      16'd489:
      begin
        register_150 <= $signed(register_150) == $signed(16'd1);
      end

      16'd490:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 567;
      end

      16'd491:
      begin
        register_150 <= 16'd7;
      end

      16'd492:
      begin
        register_150 <= $signed(register_150) + $signed(register_66);
      end

      16'd493:
      begin
        address <= register_150;
      end

      16'd494:
      begin
        register_150 <= data_out;
      end

      16'd495:
      begin
        register_150 <= data_out;
      end

      16'd496:
      begin
        register_150 <= $signed(register_150) >>> $signed(16'd8);
      end

      16'd497:
      begin
        register_150 <= $signed(register_150) & $signed(16'd15);
      end

      16'd498:
      begin
        register_150 <= $signed(register_150) << $signed(16'd1);
      end

      16'd499:
      begin
        register_69 <= register_150;
      end

      16'd500:
      begin
        register_150 <= register_69;
        register_151 <= register_69;
      end

      16'd501:
      begin
        register_150 <= $signed(register_150) + $signed(16'd7);
      end

      16'd502:
      begin
        register_70 <= register_150;
        register_150 <= 16'd8;
      end

      16'd503:
      begin
        register_150 <= $signed(register_150) + $signed(register_66);
      end

      16'd504:
      begin
        address <= register_150;
      end

      16'd505:
      begin
        register_150 <= data_out;
      end

      16'd506:
      begin
        register_150 <= data_out;
      end

      16'd507:
      begin
        register_68 <= register_150;
      end

      16'd508:
      begin
        register_150 <= register_68;
      end

      16'd509:
      begin
        register_150 <= $signed(register_150) + $signed(16'd1);
      end

      16'd510:
      begin
        register_150 <= $signed(register_150) >>> $signed(16'd1);
      end

      16'd511:
      begin
        register_150 <= $signed(register_150) - $signed(register_151);
      end

      16'd512:
      begin
        register_71 <= register_150;
        register_150 <= register_70;
      end

      16'd513:
      begin
        register_151 <= register_71;
      end

      16'd514:
      begin
        register_150 <= $signed(register_150) + $signed(register_151);
      end

      16'd515:
      begin
        register_150 <= $signed(register_150) - $signed(16'd1);
      end

      16'd516:
      begin
        register_75 <= register_150;
        register_150 <= register_70;
      end

      16'd517:
      begin
        register_150 <= $signed(register_150) + $signed(register_66);
      end

      16'd518:
      begin
        address <= register_150;
      end

      16'd519:
      begin
        register_150 <= data_out;
      end

      16'd520:
      begin
        register_150 <= data_out;
      end

      16'd521:
      begin
        register_150 <= $signed(register_150) == $signed(16'd2048);
      end

      16'd522:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 566;
      end

      16'd523:
      begin
        register_150 <= 16'd19;
      end

      16'd524:
      begin
        register_74 <= register_150;
        register_150 <= register_71;
      end

      16'd525:
      begin
        s_output_checksum <= register_150;
        program_counter <= 525;
        s_output_checksum_stb <= 1'b1;
        if (s_output_checksum_stb == 1'b1 && output_checksum_ack == 1'b1) begin
          s_output_checksum_stb <= 1'b0;
          program_counter <= 526;
        end
      end

      16'd526:
      begin
        register_150 <= 16'd0;
      end

      16'd527:
      begin
        s_output_checksum <= register_150;
        program_counter <= 527;
        s_output_checksum_stb <= 1'b1;
        if (s_output_checksum_stb == 1'b1 && output_checksum_ack == 1'b1) begin
          s_output_checksum_stb <= 1'b0;
          program_counter <= 528;
        end
      end

      16'd528:
      begin
        register_150 <= 16'd0;
      end

      16'd529:
      begin
        s_output_checksum <= register_150;
        program_counter <= 529;
        s_output_checksum_stb <= 1'b1;
        if (s_output_checksum_stb == 1'b1 && output_checksum_ack == 1'b1) begin
          s_output_checksum_stb <= 1'b0;
          program_counter <= 530;
        end
      end

      16'd530:
      begin
        register_150 <= register_70;
      end

      16'd531:
      begin
        register_150 <= $signed(register_150) + $signed(16'd2);
      end

      16'd532:
      begin
        register_73 <= register_150;
      end

      16'd533:
      begin
        register_150 <= register_73;
        register_151 <= register_75;
      end

      16'd534:
      begin
        register_150 <= $signed(register_150) <= $signed(register_151);
      end

      16'd535:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 552;
      end

      16'd536:
      begin
        register_150 <= register_73;
      end

      16'd537:
      begin
        register_150 <= $signed(register_150) + $signed(register_66);
      end

      16'd538:
      begin
        address <= register_150;
      end

      16'd539:
      begin
        register_150 <= data_out;
      end

      16'd540:
      begin
        register_150 <= data_out;
      end

      16'd541:
      begin
        register_72 <= register_150;
      end

      16'd542:
      begin
        register_150 <= register_72;
      end

      16'd543:
      begin
        s_output_checksum <= register_150;
        program_counter <= 543;
        s_output_checksum_stb <= 1'b1;
        if (s_output_checksum_stb == 1'b1 && output_checksum_ack == 1'b1) begin
          s_output_checksum_stb <= 1'b0;
          program_counter <= 544;
        end
      end

      16'd544:
      begin
        register_150 <= register_72;
        register_151 <= register_74;
      end

      16'd545:
      begin
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd546:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_74;
      end

      16'd547:
      begin
        register_150 <= $signed(register_150) + $signed(16'd1);
      end

      16'd548:
      begin
        register_74 <= register_150;
      end

      16'd549:
      begin
        register_150 <= register_73;
      end

      16'd550:
      begin
        register_150 <= $signed(register_150) + $signed(16'd1);
      end

      16'd551:
      begin
        register_73 <= register_150;
        program_counter <= 16'd533;
      end

      16'd552:
      begin
        register_150 <= 16'd0;
        register_151 <= 16'd17;
      end

      16'd553:
      begin
        register_151 <= $signed(register_151) + $signed(register_6);
      end

      16'd554:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
      end

      16'd555:
      begin
        register_150 <= input_checksum;
        program_counter <= 555;
        s_input_checksum_ack <= 1'b1;
       if (s_input_checksum_ack == 1'b1 && input_checksum_stb == 1'b1) begin
          s_input_checksum_ack <= 1'b0;
          program_counter <= 16'd556;
        end
      end

      16'd556:
      begin
        register_151 <= 16'd18;
        register_56 <= register_6;
        register_57 <= register_68;
        register_58 <= 16'd1;
        register_59 <= 16'd13;
        register_60 <= 16'd14;
      end

      16'd557:
      begin
        register_151 <= $signed(register_151) + $signed(register_6);
        register_59 <= $signed(register_59) + $signed(register_66);
        register_60 <= $signed(register_60) + $signed(register_66);
      end

      16'd558:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
      end

      16'd559:
      begin
        address <= register_59;
      end

      16'd560:
      begin
        register_59 <= data_out;
      end

      16'd561:
      begin
        register_59 <= data_out;
      end

      16'd562:
      begin
        address <= register_60;
      end

      16'd563:
      begin
        register_60 <= data_out;
      end

      16'd564:
      begin
        register_60 <= data_out;
        program_counter <= 16'd396;
        register_54 <= 16'd565;
      end

      16'd565:
      begin
        register_150 <= register_55;
        program_counter <= 16'd566;
      end

      16'd566:
      begin
        program_counter <= 16'd577;
      end

      16'd567:
      begin
        register_150 <= 16'd11;
      end

      16'd568:
      begin
        register_150 <= $signed(register_150) + $signed(register_66);
      end

      16'd569:
      begin
        address <= register_150;
      end

      16'd570:
      begin
        register_150 <= data_out;
      end

      16'd571:
      begin
        register_150 <= data_out;
      end

      16'd572:
      begin
        register_150 <= $signed(register_150) & $signed(16'd255);
      end

      16'd573:
      begin
        register_150 <= $signed(register_150) == $signed(16'd6);
      end

      16'd574:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 577;
      end

      16'd575:
      begin
        register_65 <= register_61;
        program_counter <= register_64;
      end

      16'd576:
      begin
        program_counter <= 16'd577;
      end

      16'd577:
      begin
        program_counter <= 16'd578;
      end

      16'd578:
      begin
        program_counter <= 16'd456;
      end

      16'd579:
      begin
        register_105 <= 16'd17;
        register_106 <= 16'd0;
        register_107 <= 16'd0;
        register_150 <= register_78;
      end

      16'd580:
      begin
        register_151 <= register_105;
      end

      16'd581:
      begin
        register_151 <= $signed(register_151) + $signed(16'd0);
      end

      16'd582:
      begin
        register_151 <= $signed(register_151) + $signed(register_103);
      end

      16'd583:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_79;
        register_151 <= register_105;
      end

      16'd584:
      begin
        register_151 <= $signed(register_151) + $signed(16'd1);
      end

      16'd585:
      begin
        register_151 <= $signed(register_151) + $signed(register_103);
      end

      16'd586:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd1;
        register_151 <= register_105;
      end

      16'd587:
      begin
        register_150 <= $signed(register_150) + $signed(register_80);
        register_151 <= $signed(register_151) + $signed(16'd2);
      end

      16'd588:
      begin
        address <= register_150;
        register_151 <= $signed(register_151) + $signed(register_103);
      end

      16'd589:
      begin
        register_150 <= data_out;
      end

      16'd590:
      begin
        register_150 <= data_out;
      end

      16'd591:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd0;
        register_151 <= register_105;
      end

      16'd592:
      begin
        register_150 <= $signed(register_150) + $signed(register_80);
        register_151 <= $signed(register_151) + $signed(16'd3);
      end

      16'd593:
      begin
        address <= register_150;
        register_151 <= $signed(register_151) + $signed(register_103);
      end

      16'd594:
      begin
        register_150 <= data_out;
      end

      16'd595:
      begin
        register_150 <= data_out;
      end

      16'd596:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd1;
        register_151 <= register_105;
      end

      16'd597:
      begin
        register_150 <= $signed(register_150) + $signed(register_82);
        register_151 <= $signed(register_151) + $signed(16'd4);
      end

      16'd598:
      begin
        address <= register_150;
        register_151 <= $signed(register_151) + $signed(register_103);
      end

      16'd599:
      begin
        register_150 <= data_out;
      end

      16'd600:
      begin
        register_150 <= data_out;
      end

      16'd601:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd0;
        register_151 <= register_105;
      end

      16'd602:
      begin
        register_150 <= $signed(register_150) + $signed(register_82);
        register_151 <= $signed(register_151) + $signed(16'd5);
      end

      16'd603:
      begin
        address <= register_150;
        register_151 <= $signed(register_151) + $signed(register_103);
      end

      16'd604:
      begin
        register_150 <= data_out;
      end

      16'd605:
      begin
        register_150 <= data_out;
      end

      16'd606:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd20480;
        register_151 <= register_105;
      end

      16'd607:
      begin
        register_151 <= $signed(register_151) + $signed(16'd6);
      end

      16'd608:
      begin
        register_151 <= $signed(register_151) + $signed(register_103);
      end

      16'd609:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_83;
        register_151 <= register_105;
      end

      16'd610:
      begin
        register_151 <= $signed(register_151) + $signed(16'd7);
      end

      16'd611:
      begin
        register_151 <= $signed(register_151) + $signed(register_103);
      end

      16'd612:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd0;
        register_151 <= register_105;
      end

      16'd613:
      begin
        register_151 <= $signed(register_151) + $signed(16'd8);
      end

      16'd614:
      begin
        register_151 <= $signed(register_151) + $signed(register_103);
      end

      16'd615:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd0;
        register_151 <= register_105;
      end

      16'd616:
      begin
        register_151 <= $signed(register_151) + $signed(16'd9);
      end

      16'd617:
      begin
        register_151 <= $signed(register_151) + $signed(register_103);
      end

      16'd618:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_84;
      end

      16'd619:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 628;
      end

      16'd620:
      begin
        register_150 <= register_105;
        register_151 <= register_105;
      end

      16'd621:
      begin
        register_150 <= $signed(register_150) + $signed(16'd6);
        register_151 <= $signed(register_151) + $signed(16'd6);
      end

      16'd622:
      begin
        register_150 <= $signed(register_150) + $signed(register_103);
        register_151 <= $signed(register_151) + $signed(register_103);
      end

      16'd623:
      begin
        address <= register_150;
      end

      16'd624:
      begin
        register_150 <= data_out;
      end

      16'd625:
      begin
        register_150 <= data_out;
      end

      16'd626:
      begin
        register_150 <= $signed(register_150) | $signed(16'd1);
      end

      16'd627:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        program_counter <= 16'd628;
      end

      16'd628:
      begin
        register_150 <= register_85;
      end

      16'd629:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 638;
      end

      16'd630:
      begin
        register_150 <= register_105;
        register_151 <= register_105;
      end

      16'd631:
      begin
        register_150 <= $signed(register_150) + $signed(16'd6);
        register_151 <= $signed(register_151) + $signed(16'd6);
      end

      16'd632:
      begin
        register_150 <= $signed(register_150) + $signed(register_103);
        register_151 <= $signed(register_151) + $signed(register_103);
      end

      16'd633:
      begin
        address <= register_150;
      end

      16'd634:
      begin
        register_150 <= data_out;
      end

      16'd635:
      begin
        register_150 <= data_out;
      end

      16'd636:
      begin
        register_150 <= $signed(register_150) | $signed(16'd2);
      end

      16'd637:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        program_counter <= 16'd638;
      end

      16'd638:
      begin
        register_150 <= register_86;
      end

      16'd639:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 648;
      end

      16'd640:
      begin
        register_150 <= register_105;
        register_151 <= register_105;
      end

      16'd641:
      begin
        register_150 <= $signed(register_150) + $signed(16'd6);
        register_151 <= $signed(register_151) + $signed(16'd6);
      end

      16'd642:
      begin
        register_150 <= $signed(register_150) + $signed(register_103);
        register_151 <= $signed(register_151) + $signed(register_103);
      end

      16'd643:
      begin
        address <= register_150;
      end

      16'd644:
      begin
        register_150 <= data_out;
      end

      16'd645:
      begin
        register_150 <= data_out;
      end

      16'd646:
      begin
        register_150 <= $signed(register_150) | $signed(16'd4);
      end

      16'd647:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        program_counter <= 16'd648;
      end

      16'd648:
      begin
        register_150 <= register_87;
      end

      16'd649:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 658;
      end

      16'd650:
      begin
        register_150 <= register_105;
        register_151 <= register_105;
      end

      16'd651:
      begin
        register_150 <= $signed(register_150) + $signed(16'd6);
        register_151 <= $signed(register_151) + $signed(16'd6);
      end

      16'd652:
      begin
        register_150 <= $signed(register_150) + $signed(register_103);
        register_151 <= $signed(register_151) + $signed(register_103);
      end

      16'd653:
      begin
        address <= register_150;
      end

      16'd654:
      begin
        register_150 <= data_out;
      end

      16'd655:
      begin
        register_150 <= data_out;
      end

      16'd656:
      begin
        register_150 <= $signed(register_150) | $signed(16'd8);
      end

      16'd657:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        program_counter <= 16'd658;
      end

      16'd658:
      begin
        register_150 <= register_88;
      end

      16'd659:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 668;
      end

      16'd660:
      begin
        register_150 <= register_105;
        register_151 <= register_105;
      end

      16'd661:
      begin
        register_150 <= $signed(register_150) + $signed(16'd6);
        register_151 <= $signed(register_151) + $signed(16'd6);
      end

      16'd662:
      begin
        register_150 <= $signed(register_150) + $signed(register_103);
        register_151 <= $signed(register_151) + $signed(register_103);
      end

      16'd663:
      begin
        address <= register_150;
      end

      16'd664:
      begin
        register_150 <= data_out;
      end

      16'd665:
      begin
        register_150 <= data_out;
      end

      16'd666:
      begin
        register_150 <= $signed(register_150) | $signed(16'd16);
      end

      16'd667:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        program_counter <= 16'd668;
      end

      16'd668:
      begin
        register_150 <= register_89;
      end

      16'd669:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 678;
      end

      16'd670:
      begin
        register_150 <= register_105;
        register_151 <= register_105;
      end

      16'd671:
      begin
        register_150 <= $signed(register_150) + $signed(16'd6);
        register_151 <= $signed(register_151) + $signed(16'd6);
      end

      16'd672:
      begin
        register_150 <= $signed(register_150) + $signed(register_103);
        register_151 <= $signed(register_151) + $signed(register_103);
      end

      16'd673:
      begin
        address <= register_150;
      end

      16'd674:
      begin
        register_150 <= data_out;
      end

      16'd675:
      begin
        register_150 <= data_out;
      end

      16'd676:
      begin
        register_150 <= $signed(register_150) | $signed(16'd32);
      end

      16'd677:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        program_counter <= 16'd678;
      end

      16'd678:
      begin
        program_counter <= 16'd2;
        register_8 <= 16'd679;
      end

      16'd679:
      begin
        register_150 <= register_9;
        register_12 <= register_3;
        program_counter <= 16'd7;
        register_10 <= 16'd680;
      end

      16'd680:
      begin
        register_150 <= register_11;
        register_12 <= register_4;
        program_counter <= 16'd7;
        register_10 <= 16'd681;
      end

      16'd681:
      begin
        register_150 <= register_11;
        register_12 <= register_76;
        program_counter <= 16'd7;
        register_10 <= 16'd682;
      end

      16'd682:
      begin
        register_150 <= register_11;
        register_12 <= register_77;
        program_counter <= 16'd7;
        register_10 <= 16'd683;
      end

      16'd683:
      begin
        register_150 <= register_11;
        register_12 <= 16'd6;
        program_counter <= 16'd7;
        register_10 <= 16'd684;
      end

      16'd684:
      begin
        register_150 <= register_11;
        register_12 <= register_104;
      end

      16'd685:
      begin
        register_12 <= $signed(register_12) + $signed(16'd20);
        program_counter <= 16'd7;
        register_10 <= 16'd686;
      end

      16'd686:
      begin
        register_150 <= register_11;
      end

      16'd687:
      begin
        register_150 <= register_104;
      end

      16'd688:
      begin
        register_150 <= $signed(register_150) + $signed(16'd20);
      end

      16'd689:
      begin
        register_150 <= $signed(register_150) + $signed(16'd1);
      end

      16'd690:
      begin
        register_150 <= $signed(register_150) >>> $signed(16'd1);
      end

      16'd691:
      begin
        register_106 <= register_150;
        register_150 <= register_105;
      end

      16'd692:
      begin
        register_107 <= register_150;
        register_150 <= 16'd0;
      end

      16'd693:
      begin
        register_72 <= register_150;
      end

      16'd694:
      begin
        register_150 <= register_72;
        register_151 <= register_106;
      end

      16'd695:
      begin
        register_150 <= $signed(register_150) < $signed(register_151);
      end

      16'd696:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 709;
      end

      16'd697:
      begin
        register_12 <= register_107;
      end

      16'd698:
      begin
        register_12 <= $signed(register_12) + $signed(register_103);
      end

      16'd699:
      begin
        address <= register_12;
      end

      16'd700:
      begin
        register_12 <= data_out;
      end

      16'd701:
      begin
        register_12 <= data_out;
        program_counter <= 16'd7;
        register_10 <= 16'd702;
      end

      16'd702:
      begin
        register_150 <= register_11;
      end

      16'd703:
      begin
        register_150 <= register_107;
      end

      16'd704:
      begin
        register_150 <= $signed(register_150) + $signed(16'd1);
      end

      16'd705:
      begin
        register_107 <= register_150;
      end

      16'd706:
      begin
        register_150 <= register_72;
      end

      16'd707:
      begin
        register_150 <= $signed(register_150) + $signed(16'd1);
      end

      16'd708:
      begin
        register_72 <= register_150;
        program_counter <= 16'd694;
      end

      16'd709:
      begin
        program_counter <= 16'd36;
        register_14 <= 16'd710;
      end

      16'd710:
      begin
        register_150 <= register_15;
        register_151 <= register_105;
        register_56 <= register_103;
        register_57 <= register_104;
        register_58 <= 16'd6;
        register_59 <= register_76;
        register_60 <= register_77;
      end

      16'd711:
      begin
        register_151 <= $signed(register_151) + $signed(16'd8);
        register_57 <= $signed(register_57) + $signed(16'd40);
      end

      16'd712:
      begin
        register_151 <= $signed(register_151) + $signed(register_103);
      end

      16'd713:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        program_counter <= 16'd396;
        register_54 <= 16'd714;
      end

      16'd714:
      begin
        register_150 <= register_55;
        register_102 <= 16'd0;
        program_counter <= register_101;
      end

      16'd715:
      begin
        register_113 <= 16'd0;
        register_114 <= 16'd0;
        register_115 <= 16'd0;
        register_116 <= 16'd0;
        register_117 <= 16'd0;
        register_118 <= 16'd0;
        register_119 <= 16'd0;
        register_66 <= register_112;
        program_counter <= 16'd455;
        register_64 <= 16'd716;
      end

      16'd716:
      begin
        register_150 <= register_65;
        register_111 <= 16'd0;
      end

      16'd717:
      begin
        register_113 <= register_150;
        register_150 <= 16'd7;
      end

      16'd718:
      begin
        register_150 <= $signed(register_150) + $signed(register_112);
      end

      16'd719:
      begin
        address <= register_150;
      end

      16'd720:
      begin
        register_150 <= data_out;
      end

      16'd721:
      begin
        register_150 <= data_out;
      end

      16'd722:
      begin
        register_150 <= $signed(register_150) >>> $signed(16'd8);
      end

      16'd723:
      begin
        register_150 <= $signed(register_150) & $signed(16'd15);
      end

      16'd724:
      begin
        register_150 <= $signed(register_150) << $signed(16'd1);
      end

      16'd725:
      begin
        register_114 <= register_150;
      end

      16'd726:
      begin
        register_150 <= register_114;
        register_151 <= register_114;
      end

      16'd727:
      begin
        register_150 <= $signed(register_150) + $signed(16'd7);
        register_151 <= $signed(register_151) << $signed(16'd1);
      end

      16'd728:
      begin
        register_115 <= register_150;
        register_150 <= 16'd8;
      end

      16'd729:
      begin
        register_150 <= $signed(register_150) + $signed(register_112);
      end

      16'd730:
      begin
        address <= register_150;
      end

      16'd731:
      begin
        register_150 <= data_out;
      end

      16'd732:
      begin
        register_150 <= data_out;
      end

      16'd733:
      begin
        register_116 <= register_150;
      end

      16'd734:
      begin
        register_150 <= register_116;
      end

      16'd735:
      begin
        register_150 <= $signed(register_150) - $signed(register_151);
      end

      16'd736:
      begin
        register_117 <= register_150;
        register_150 <= register_115;
      end

      16'd737:
      begin
        register_150 <= $signed(register_150) + $signed(16'd6);
      end

      16'd738:
      begin
        register_150 <= $signed(register_150) + $signed(register_112);
      end

      16'd739:
      begin
        address <= register_150;
      end

      16'd740:
      begin
        register_150 <= data_out;
      end

      16'd741:
      begin
        register_150 <= data_out;
      end

      16'd742:
      begin
        register_150 <= $signed(register_150) & $signed(16'd61440);
      end

      16'd743:
      begin
        register_150 <= $signed(register_150) >>> $signed(16'd10);
      end

      16'd744:
      begin
        register_119 <= register_150;
        register_150 <= register_117;
      end

      16'd745:
      begin
        register_151 <= register_119;
      end

      16'd746:
      begin
        register_150 <= $signed(register_150) - $signed(register_151);
        register_151 <= register_119;
      end

      16'd747:
      begin
        register_108 <= register_150;
        register_150 <= register_115;
        register_151 <= $signed(register_151) >>> $signed(16'd1);
      end

      16'd748:
      begin
        register_150 <= $signed(register_150) + $signed(register_151);
        register_151 <= 16'd1;
      end

      16'd749:
      begin
        register_109 <= register_150;
        register_150 <= register_115;
        register_151 <= $signed(register_151) + $signed(register_92);
      end

      16'd750:
      begin
        register_150 <= $signed(register_150) + $signed(16'd0);
      end

      16'd751:
      begin
        register_150 <= $signed(register_150) + $signed(register_112);
      end

      16'd752:
      begin
        address <= register_150;
      end

      16'd753:
      begin
        register_150 <= data_out;
      end

      16'd754:
      begin
        register_150 <= data_out;
      end

      16'd755:
      begin
        register_90 <= register_150;
        register_150 <= register_115;
      end

      16'd756:
      begin
        register_150 <= $signed(register_150) + $signed(16'd1);
      end

      16'd757:
      begin
        register_150 <= $signed(register_150) + $signed(register_112);
      end

      16'd758:
      begin
        address <= register_150;
      end

      16'd759:
      begin
        register_150 <= data_out;
      end

      16'd760:
      begin
        register_150 <= data_out;
      end

      16'd761:
      begin
        register_91 <= register_150;
        register_150 <= register_115;
      end

      16'd762:
      begin
        register_150 <= $signed(register_150) + $signed(16'd2);
      end

      16'd763:
      begin
        register_150 <= $signed(register_150) + $signed(register_112);
      end

      16'd764:
      begin
        address <= register_150;
      end

      16'd765:
      begin
        register_150 <= data_out;
      end

      16'd766:
      begin
        register_150 <= data_out;
      end

      16'd767:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_115;
        register_151 <= 16'd0;
      end

      16'd768:
      begin
        register_150 <= $signed(register_150) + $signed(16'd3);
        register_151 <= $signed(register_151) + $signed(register_92);
      end

      16'd769:
      begin
        register_150 <= $signed(register_150) + $signed(register_112);
      end

      16'd770:
      begin
        address <= register_150;
      end

      16'd771:
      begin
        register_150 <= data_out;
      end

      16'd772:
      begin
        register_150 <= data_out;
      end

      16'd773:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_115;
        register_151 <= 16'd1;
      end

      16'd774:
      begin
        register_150 <= $signed(register_150) + $signed(16'd4);
        register_151 <= $signed(register_151) + $signed(register_93);
      end

      16'd775:
      begin
        register_150 <= $signed(register_150) + $signed(register_112);
      end

      16'd776:
      begin
        address <= register_150;
      end

      16'd777:
      begin
        register_150 <= data_out;
      end

      16'd778:
      begin
        register_150 <= data_out;
      end

      16'd779:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_115;
        register_151 <= 16'd0;
      end

      16'd780:
      begin
        register_150 <= $signed(register_150) + $signed(16'd5);
        register_151 <= $signed(register_151) + $signed(register_93);
      end

      16'd781:
      begin
        register_150 <= $signed(register_150) + $signed(register_112);
      end

      16'd782:
      begin
        address <= register_150;
      end

      16'd783:
      begin
        register_150 <= data_out;
      end

      16'd784:
      begin
        register_150 <= data_out;
      end

      16'd785:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_115;
      end

      16'd786:
      begin
        register_150 <= $signed(register_150) + $signed(16'd7);
      end

      16'd787:
      begin
        register_150 <= $signed(register_150) + $signed(register_112);
      end

      16'd788:
      begin
        address <= register_150;
      end

      16'd789:
      begin
        register_150 <= data_out;
      end

      16'd790:
      begin
        register_150 <= data_out;
      end

      16'd791:
      begin
        register_94 <= register_150;
        register_150 <= register_115;
      end

      16'd792:
      begin
        register_150 <= $signed(register_150) + $signed(16'd6);
      end

      16'd793:
      begin
        register_150 <= $signed(register_150) + $signed(register_112);
      end

      16'd794:
      begin
        address <= register_150;
      end

      16'd795:
      begin
        register_150 <= data_out;
      end

      16'd796:
      begin
        register_150 <= data_out;
      end

      16'd797:
      begin
        register_150 <= $signed(register_150) & $signed(16'd1);
      end

      16'd798:
      begin
        register_95 <= register_150;
        register_150 <= register_115;
      end

      16'd799:
      begin
        register_150 <= $signed(register_150) + $signed(16'd6);
      end

      16'd800:
      begin
        register_150 <= $signed(register_150) + $signed(register_112);
      end

      16'd801:
      begin
        address <= register_150;
      end

      16'd802:
      begin
        register_150 <= data_out;
      end

      16'd803:
      begin
        register_150 <= data_out;
      end

      16'd804:
      begin
        register_150 <= $signed(register_150) & $signed(16'd2);
      end

      16'd805:
      begin
        register_96 <= register_150;
        register_150 <= register_115;
      end

      16'd806:
      begin
        register_150 <= $signed(register_150) + $signed(16'd6);
      end

      16'd807:
      begin
        register_150 <= $signed(register_150) + $signed(register_112);
      end

      16'd808:
      begin
        address <= register_150;
      end

      16'd809:
      begin
        register_150 <= data_out;
      end

      16'd810:
      begin
        register_150 <= data_out;
      end

      16'd811:
      begin
        register_150 <= $signed(register_150) & $signed(16'd4);
      end

      16'd812:
      begin
        register_97 <= register_150;
        register_150 <= register_115;
      end

      16'd813:
      begin
        register_150 <= $signed(register_150) + $signed(16'd6);
      end

      16'd814:
      begin
        register_150 <= $signed(register_150) + $signed(register_112);
      end

      16'd815:
      begin
        address <= register_150;
      end

      16'd816:
      begin
        register_150 <= data_out;
      end

      16'd817:
      begin
        register_150 <= data_out;
      end

      16'd818:
      begin
        register_150 <= $signed(register_150) & $signed(16'd8);
      end

      16'd819:
      begin
        register_98 <= register_150;
        register_150 <= register_115;
      end

      16'd820:
      begin
        register_150 <= $signed(register_150) + $signed(16'd6);
      end

      16'd821:
      begin
        register_150 <= $signed(register_150) + $signed(register_112);
      end

      16'd822:
      begin
        address <= register_150;
      end

      16'd823:
      begin
        register_150 <= data_out;
      end

      16'd824:
      begin
        register_150 <= data_out;
      end

      16'd825:
      begin
        register_150 <= $signed(register_150) & $signed(16'd16);
      end

      16'd826:
      begin
        register_99 <= register_150;
        register_150 <= register_115;
      end

      16'd827:
      begin
        register_150 <= $signed(register_150) + $signed(16'd6);
      end

      16'd828:
      begin
        register_150 <= $signed(register_150) + $signed(register_112);
      end

      16'd829:
      begin
        address <= register_150;
      end

      16'd830:
      begin
        register_150 <= data_out;
      end

      16'd831:
      begin
        register_150 <= data_out;
      end

      16'd832:
      begin
        register_150 <= $signed(register_150) & $signed(16'd32);
      end

      16'd833:
      begin
        register_100 <= register_150;
        program_counter <= register_110;
      end

      16'd834:
      begin
        register_125 <= 16'd0;
        register_126 <= 16'd0;
        register_127 <= 16'd0;
        register_150 <= register_123;
      end

      16'd835:
      begin
        register_126 <= register_150;
        register_150 <= register_124;
      end

      16'd836:
      begin
        register_125 <= register_150;
      end

      16'd837:
      begin
        register_150 <= register_125;
      end

      16'd838:
      begin
        register_150 <= $signed(register_150) > $signed(16'd0);
      end

      16'd839:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 861;
      end

      16'd840:
      begin
        register_150 <= register_126;
      end

      16'd841:
      begin
        register_150 <= $signed(register_150) + $signed(register_122);
      end

      16'd842:
      begin
        address <= register_150;
      end

      16'd843:
      begin
        register_150 <= data_out;
      end

      16'd844:
      begin
        register_150 <= data_out;
      end

      16'd845:
      begin
        register_127 <= register_150;
        register_150 <= register_125;
      end

      16'd846:
      begin
        register_150 <= $signed(register_150) > $signed(16'd1);
      end

      16'd847:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 852;
      end

      16'd848:
      begin
        register_150 <= register_127;
      end

      16'd849:
      begin
        register_150 <= $signed(register_150) >>> $signed(16'd8);
      end

      16'd850:
      begin
        s_output_rs232_tx <= register_150;
        program_counter <= 850;
        s_output_rs232_tx_stb <= 1'b1;
        if (s_output_rs232_tx_stb == 1'b1 && output_rs232_tx_ack == 1'b1) begin
          s_output_rs232_tx_stb <= 1'b0;
          program_counter <= 851;
        end
      end

      16'd851:
      begin
        program_counter <= 16'd852;
      end

      16'd852:
      begin
        register_150 <= register_127;
      end

      16'd853:
      begin
        register_150 <= $signed(register_150) & $signed(16'd255);
      end

      16'd854:
      begin
        s_output_rs232_tx <= register_150;
        program_counter <= 854;
        s_output_rs232_tx_stb <= 1'b1;
        if (s_output_rs232_tx_stb == 1'b1 && output_rs232_tx_ack == 1'b1) begin
          s_output_rs232_tx_stb <= 1'b0;
          program_counter <= 855;
        end
      end

      16'd855:
      begin
        register_150 <= register_126;
      end

      16'd856:
      begin
        register_150 <= $signed(register_150) + $signed(16'd1);
      end

      16'd857:
      begin
        register_126 <= register_150;
      end

      16'd858:
      begin
        register_150 <= register_125;
      end

      16'd859:
      begin
        register_150 <= $signed(register_150) - $signed(16'd2);
      end

      16'd860:
      begin
        register_125 <= register_150;
        program_counter <= 16'd837;
      end

      16'd861:
      begin
        register_121 <= 16'd0;
        program_counter <= register_120;
      end

      16'd862:
      begin
        register_132 <= 16'd620;
        register_133 <= 16'd0;
        register_134 <= 16'd0;
        register_135 <= 16'd0;
        register_150 <= register_131;
      end

      16'd863:
      begin
        register_135 <= register_150;
        register_150 <= 16'd0;
      end

      16'd864:
      begin
        register_133 <= register_150;
      end

      16'd865:
      begin
        register_150 <= register_133;
      end

      16'd866:
      begin
        register_150 <= $signed(register_150) + $signed(register_132);
      end

      16'd867:
      begin
        address <= register_150;
      end

      16'd868:
      begin
        register_150 <= data_out;
      end

      16'd869:
      begin
        register_150 <= data_out;
      end

      16'd870:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 878;
      end

      16'd871:
      begin
        register_150 <= register_133;
      end

      16'd872:
      begin
        register_150 <= $signed(register_150) + $signed(register_132);
      end

      16'd873:
      begin
        address <= register_150;
      end

      16'd874:
      begin
        register_150 <= data_out;
      end

      16'd875:
      begin
        register_150 <= data_out;
      end

      16'd876:
      begin
        register_150 <= $signed(register_150) << $signed(16'd8);
      end

      16'd877:
      begin
        register_134 <= register_150;
        program_counter <= 16'd879;
      end

      16'd878:
      begin
        program_counter <= 16'd905;
      end

      16'd879:
      begin
        register_150 <= register_133;
      end

      16'd880:
      begin
        register_150 <= $signed(register_150) + $signed(16'd1);
      end

      16'd881:
      begin
        register_133 <= register_150;
      end

      16'd882:
      begin
        register_150 <= register_133;
      end

      16'd883:
      begin
        register_150 <= $signed(register_150) + $signed(register_132);
      end

      16'd884:
      begin
        address <= register_150;
      end

      16'd885:
      begin
        register_150 <= data_out;
      end

      16'd886:
      begin
        register_150 <= data_out;
      end

      16'd887:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 895;
      end

      16'd888:
      begin
        register_150 <= register_134;
        register_151 <= register_133;
      end

      16'd889:
      begin
        register_151 <= $signed(register_151) + $signed(register_132);
      end

      16'd890:
      begin
        address <= register_151;
      end

      16'd891:
      begin
        register_151 <= data_out;
      end

      16'd892:
      begin
        register_151 <= data_out;
      end

      16'd893:
      begin
        register_150 <= $signed(register_150) | $signed(register_151);
      end

      16'd894:
      begin
        register_134 <= register_150;
        program_counter <= 16'd898;
      end

      16'd895:
      begin
        register_150 <= register_134;
        register_151 <= register_135;
      end

      16'd896:
      begin
        register_151 <= $signed(register_151) + $signed(register_130);
      end

      16'd897:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        program_counter <= 16'd905;
      end

      16'd898:
      begin
        register_150 <= register_134;
        register_151 <= register_135;
      end

      16'd899:
      begin
        register_151 <= $signed(register_151) + $signed(register_130);
      end

      16'd900:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= register_133;
      end

      16'd901:
      begin
        register_150 <= $signed(register_150) + $signed(16'd1);
      end

      16'd902:
      begin
        register_133 <= register_150;
        register_150 <= register_135;
      end

      16'd903:
      begin
        register_150 <= $signed(register_150) + $signed(16'd1);
      end

      16'd904:
      begin
        register_135 <= register_150;
        program_counter <= 16'd865;
      end

      16'd905:
      begin
        register_129 <= register_133;
        program_counter <= register_128;
      end

      16'd906:
      begin
        register_138 <= 16'd646;
        register_139 <= 16'd1670;
        register_140 <= 16'd27;
        register_141 <= 16'd1;
        register_142 <= 16'd2;
        register_143 <= 16'd3;
        register_144 <= 16'd4;
        register_146 <= 16'd0;
        register_147 <= 16'd0;
        register_148 <= 16'd0;
        register_149 <= 16'd0;
        register_150 <= 16'd0;
        register_151 <= 16'd0;
      end

      16'd907:
      begin
        register_145 <= register_141;
        register_151 <= $signed(register_151) + $signed(register_80);
      end

      16'd908:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd0;
        register_151 <= 16'd1;
      end

      16'd909:
      begin
        register_151 <= $signed(register_151) + $signed(register_80);
      end

      16'd910:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
      end

      16'd911:
      begin
        register_150 <= register_145;
        register_151 <= register_141;
      end

      16'd912:
      begin
        register_150 <= $signed(register_150) == $signed(register_151);
      end

      16'd913:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 944;
      end

      16'd914:
      begin
        register_112 <= register_138;
        program_counter <= 16'd715;
        register_110 <= 16'd915;
      end

      16'd915:
      begin
        register_150 <= register_111;
        register_151 <= register_5;
      end

      16'd916:
      begin
        register_150 <= register_91;
      end

      16'd917:
      begin
        register_150 <= $signed(register_150) == $signed(register_151);
      end

      16'd918:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 921;
      end

      16'd919:
      begin
        program_counter <= 16'd922;
      end

      16'd920:
      begin
        program_counter <= 16'd921;
      end

      16'd921:
      begin
        program_counter <= 16'd914;
      end

      16'd922:
      begin
        register_150 <= register_96;
      end

      16'd923:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 943;
      end

      16'd924:
      begin
        register_150 <= 16'd13;
        register_18 <= register_82;
        register_19 <= register_92;
        register_20 <= 16'd1;
      end

      16'd925:
      begin
        register_150 <= $signed(register_150) + $signed(register_138);
      end

      16'd926:
      begin
        address <= register_150;
      end

      16'd927:
      begin
        register_150 <= data_out;
      end

      16'd928:
      begin
        register_150 <= data_out;
      end

      16'd929:
      begin
        register_76 <= register_150;
        register_150 <= 16'd14;
      end

      16'd930:
      begin
        register_150 <= $signed(register_150) + $signed(register_138);
      end

      16'd931:
      begin
        address <= register_150;
      end

      16'd932:
      begin
        register_150 <= data_out;
      end

      16'd933:
      begin
        register_150 <= data_out;
      end

      16'd934:
      begin
        register_77 <= register_150;
        register_150 <= register_90;
      end

      16'd935:
      begin
        register_79 <= register_150;
        register_150 <= register_5;
      end

      16'd936:
      begin
        register_78 <= register_150;
        program_counter <= 16'd46;
        register_16 <= 16'd937;
      end

      16'd937:
      begin
        register_150 <= register_17;
        register_103 <= register_139;
        register_104 <= 16'd0;
      end

      16'd938:
      begin
        register_150 <= 16'd1;
      end

      16'd939:
      begin
        register_85 <= register_150;
        register_150 <= 16'd1;
      end

      16'd940:
      begin
        register_88 <= register_150;
        register_150 <= register_142;
      end

      16'd941:
      begin
        register_145 <= register_150;
        program_counter <= 16'd579;
        register_101 <= 16'd942;
      end

      16'd942:
      begin
        register_150 <= register_102;
        program_counter <= 16'd943;
      end

      16'd943:
      begin
        program_counter <= 16'd1068;
      end

      16'd944:
      begin
        register_150 <= register_145;
        register_151 <= register_142;
      end

      16'd945:
      begin
        register_150 <= $signed(register_150) == $signed(register_151);
      end

      16'd946:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 982;
      end

      16'd947:
      begin
        register_112 <= register_138;
        program_counter <= 16'd715;
        register_110 <= 16'd948;
      end

      16'd948:
      begin
        register_150 <= register_111;
        register_151 <= register_5;
      end

      16'd949:
      begin
        register_150 <= register_91;
      end

      16'd950:
      begin
        register_150 <= $signed(register_150) == $signed(register_151);
      end

      16'd951:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 954;
      end

      16'd952:
      begin
        program_counter <= 16'd955;
      end

      16'd953:
      begin
        program_counter <= 16'd954;
      end

      16'd954:
      begin
        program_counter <= 16'd947;
      end

      16'd955:
      begin
        register_150 <= register_99;
      end

      16'd956:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 981;
      end

      16'd957:
      begin
        register_150 <= register_143;
        register_151 <= 16'd1;
      end

      16'd958:
      begin
        register_145 <= register_150;
        register_150 <= 16'd1;
        register_151 <= $signed(register_151) + $signed(register_80);
      end

      16'd959:
      begin
        register_150 <= $signed(register_150) + $signed(register_93);
      end

      16'd960:
      begin
        address <= register_150;
      end

      16'd961:
      begin
        register_150 <= data_out;
      end

      16'd962:
      begin
        register_150 <= data_out;
      end

      16'd963:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd0;
        register_151 <= 16'd0;
      end

      16'd964:
      begin
        register_150 <= $signed(register_150) + $signed(register_93);
        register_151 <= $signed(register_151) + $signed(register_80);
      end

      16'd965:
      begin
        address <= register_150;
      end

      16'd966:
      begin
        register_150 <= data_out;
      end

      16'd967:
      begin
        register_150 <= data_out;
      end

      16'd968:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd1;
        register_151 <= 16'd1;
      end

      16'd969:
      begin
        register_150 <= $signed(register_150) + $signed(register_93);
        register_151 <= $signed(register_151) + $signed(register_81);
      end

      16'd970:
      begin
        address <= register_150;
      end

      16'd971:
      begin
        register_150 <= data_out;
      end

      16'd972:
      begin
        register_150 <= data_out;
      end

      16'd973:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd0;
        register_151 <= 16'd0;
      end

      16'd974:
      begin
        register_150 <= $signed(register_150) + $signed(register_93);
        register_151 <= $signed(register_151) + $signed(register_81);
      end

      16'd975:
      begin
        address <= register_150;
      end

      16'd976:
      begin
        register_150 <= data_out;
      end

      16'd977:
      begin
        register_150 <= data_out;
      end

      16'd978:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd0;
      end

      16'd979:
      begin
        register_85 <= register_150;
        register_150 <= 16'd0;
      end

      16'd980:
      begin
        register_88 <= register_150;
        program_counter <= 16'd981;
      end

      16'd981:
      begin
        program_counter <= 16'd1068;
      end

      16'd982:
      begin
        register_150 <= register_145;
        register_151 <= register_143;
      end

      16'd983:
      begin
        register_150 <= $signed(register_150) == $signed(register_151);
      end

      16'd984:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 1049;
      end

      16'd985:
      begin
        register_112 <= register_138;
        program_counter <= 16'd715;
        register_110 <= 16'd986;
      end

      16'd986:
      begin
        register_150 <= register_111;
        register_151 <= register_5;
      end

      16'd987:
      begin
        register_150 <= register_91;
      end

      16'd988:
      begin
        register_150 <= $signed(register_150) == $signed(register_151);
      end

      16'd989:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 992;
      end

      16'd990:
      begin
        program_counter <= 16'd993;
      end

      16'd991:
      begin
        program_counter <= 16'd992;
      end

      16'd992:
      begin
        program_counter <= 16'd985;
      end

      16'd993:
      begin
        register_150 <= 16'd1;
      end

      16'd994:
      begin
        register_88 <= register_150;
        register_150 <= register_95;
      end

      16'd995:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 1003;
      end

      16'd996:
      begin
        register_150 <= 16'd1;
        register_18 <= register_82;
        register_19 <= register_92;
        register_20 <= 16'd1;
      end

      16'd997:
      begin
        register_88 <= register_150;
        register_150 <= 16'd1;
      end

      16'd998:
      begin
        register_84 <= register_150;
        program_counter <= 16'd46;
        register_16 <= 16'd999;
      end

      16'd999:
      begin
        register_150 <= register_17;
        register_103 <= register_139;
        register_104 <= 16'd0;
      end

      16'd1000:
      begin
        register_150 <= register_144;
      end

      16'd1001:
      begin
        register_145 <= register_150;
        program_counter <= 16'd579;
        register_101 <= 16'd1002;
      end

      16'd1002:
      begin
        register_150 <= register_102;
        program_counter <= 16'd1048;
      end

      16'd1003:
      begin
        register_18 <= register_82;
        register_19 <= register_92;
        register_20 <= register_108;
        program_counter <= 16'd46;
        register_16 <= 16'd1004;
      end

      16'd1004:
      begin
        register_150 <= register_17;
      end

      16'd1005:
      begin
        register_146 <= register_150;
      end

      16'd1006:
      begin
        register_150 <= register_146;
      end

      16'd1007:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 1010;
      end

      16'd1008:
      begin
        register_122 <= register_138;
        register_123 <= register_109;
        register_124 <= register_108;
        program_counter <= 16'd834;
        register_120 <= 16'd1009;
      end

      16'd1009:
      begin
        register_150 <= register_121;
        program_counter <= 16'd1010;
      end

      16'd1010:
      begin
        register_150 <= register_99;
      end

      16'd1011:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 1021;
      end

      16'd1012:
      begin
        register_150 <= 16'd1;
        register_151 <= 16'd1;
      end

      16'd1013:
      begin
        register_150 <= $signed(register_150) + $signed(register_81);
        register_151 <= $signed(register_151) + $signed(register_93);
      end

      16'd1014:
      begin
        address <= register_150;
      end

      16'd1015:
      begin
        register_150 <= data_out;
      end

      16'd1016:
      begin
        register_150 <= data_out;
      end

      16'd1017:
      begin
        address <= register_151;
      end

      16'd1018:
      begin
        register_151 <= data_out;
      end

      16'd1019:
      begin
        register_151 <= data_out;
      end

      16'd1020:
      begin
        register_150 <= $signed(register_150) == $signed(register_151);
      end

      16'd1021:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 1031;
      end

      16'd1022:
      begin
        register_150 <= 16'd0;
        register_151 <= 16'd0;
      end

      16'd1023:
      begin
        register_150 <= $signed(register_150) + $signed(register_81);
        register_151 <= $signed(register_151) + $signed(register_93);
      end

      16'd1024:
      begin
        address <= register_150;
      end

      16'd1025:
      begin
        register_150 <= data_out;
      end

      16'd1026:
      begin
        register_150 <= data_out;
      end

      16'd1027:
      begin
        address <= register_151;
      end

      16'd1028:
      begin
        register_151 <= data_out;
      end

      16'd1029:
      begin
        register_151 <= data_out;
      end

      16'd1030:
      begin
        register_150 <= $signed(register_150) == $signed(register_151);
      end

      16'd1031:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 1046;
      end

      16'd1032:
      begin
        register_130 <= register_139;
        register_131 <= register_140;
        program_counter <= 16'd862;
        register_128 <= 16'd1033;
      end

      16'd1033:
      begin
        register_150 <= register_129;
        register_151 <= 16'd0;
        register_18 <= register_81;
        register_19 <= register_80;
      end

      16'd1034:
      begin
        register_148 <= register_150;
        register_150 <= 16'd0;
        register_151 <= $signed(register_151) + $signed(register_80);
      end

      16'd1035:
      begin
        register_150 <= $signed(register_150) + $signed(register_81);
        register_20 <= register_148;
      end

      16'd1036:
      begin
        address <= register_150;
      end

      16'd1037:
      begin
        register_150 <= data_out;
      end

      16'd1038:
      begin
        register_150 <= data_out;
      end

      16'd1039:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        register_150 <= 16'd1;
        register_151 <= 16'd1;
      end

      16'd1040:
      begin
        register_150 <= $signed(register_150) + $signed(register_81);
        register_151 <= $signed(register_151) + $signed(register_80);
      end

      16'd1041:
      begin
        address <= register_150;
      end

      16'd1042:
      begin
        register_150 <= data_out;
      end

      16'd1043:
      begin
        register_150 <= data_out;
      end

      16'd1044:
      begin
        address <= register_151;
        data_in <= register_150;
        write_enable <= 1'b1;
        program_counter <= 16'd46;
        register_16 <= 16'd1045;
      end

      16'd1045:
      begin
        register_150 <= register_17;
        program_counter <= 16'd1046;
      end

      16'd1046:
      begin
        register_103 <= register_139;
        register_104 <= register_148;
        program_counter <= 16'd579;
        register_101 <= 16'd1047;
      end

      16'd1047:
      begin
        register_150 <= register_102;
      end

      16'd1048:
      begin
        program_counter <= 16'd1068;
      end

      16'd1049:
      begin
        register_150 <= register_145;
        register_151 <= register_144;
      end

      16'd1050:
      begin
        register_150 <= $signed(register_150) == $signed(register_151);
      end

      16'd1051:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 1068;
      end

      16'd1052:
      begin
        register_112 <= register_138;
        program_counter <= 16'd715;
        register_110 <= 16'd1053;
      end

      16'd1053:
      begin
        register_150 <= register_111;
        register_151 <= register_5;
      end

      16'd1054:
      begin
        register_150 <= register_91;
      end

      16'd1055:
      begin
        register_150 <= $signed(register_150) == $signed(register_151);
      end

      16'd1056:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 1059;
      end

      16'd1057:
      begin
        program_counter <= 16'd1060;
      end

      16'd1058:
      begin
        program_counter <= 16'd1059;
      end

      16'd1059:
      begin
        program_counter <= 16'd1052;
      end

      16'd1060:
      begin
        register_150 <= register_99;
      end

      16'd1061:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 1067;
      end

      16'd1062:
      begin
        register_150 <= register_141;
      end

      16'd1063:
      begin
        register_145 <= register_150;
        register_150 <= 16'd0;
      end

      16'd1064:
      begin
        register_85 <= register_150;
        register_150 <= 16'd0;
      end

      16'd1065:
      begin
        register_84 <= register_150;
        register_150 <= 16'd0;
      end

      16'd1066:
      begin
        register_88 <= register_150;
        program_counter <= 16'd1067;
      end

      16'd1067:
      begin
        program_counter <= 16'd1068;
      end

      16'd1068:
      begin
        register_150 <= register_97;
      end

      16'd1069:
      begin
        if (register_150 == 16'h0000)
          program_counter <= 1072;
      end

      16'd1070:
      begin
        register_150 <= register_141;
      end

      16'd1071:
      begin
        register_145 <= register_150;
        program_counter <= 16'd1072;
      end

      16'd1072:
      begin
        program_counter <= 16'd911;
      end

      16'd1073:
      begin
        register_150 <= 16'd5;
      end

      16'd1074:
      begin
        s_output_leds <= register_150;
        program_counter <= 1074;
        s_output_leds_stb <= 1'b1;
        if (s_output_leds_stb == 1'b1 && output_leds_ack == 1'b1) begin
          s_output_leds_stb <= 1'b0;
          program_counter <= 1075;
        end
      end

      16'd1075:
      begin
        register_150 <= input_rs232_rx;
        program_counter <= 1075;
        s_input_rs232_rx_ack <= 1'b1;
       if (s_input_rs232_rx_ack == 1'b1 && input_rs232_rx_stb == 1'b1) begin
          s_input_rs232_rx_ack <= 1'b0;
          program_counter <= 16'd1076;
        end
      end

      16'd1076:
      begin
        register_150 <= 16'd1;
      end

      16'd1077:
      begin
        s_output_rs232_tx <= register_150;
        program_counter <= 1077;
        s_output_rs232_tx_stb <= 1'b1;
        if (s_output_rs232_tx_stb == 1'b1 && output_rs232_tx_ack == 1'b1) begin
          s_output_rs232_tx_stb <= 1'b0;
          program_counter <= 1078;
        end
      end

      16'd1078:
      begin
        register_137 <= 16'd0;
        program_counter <= register_136;
      end

    endcase
    if (rst == 1'b1) begin
      program_counter <= 0;
    end
  end
  assign input_checksum_ack = s_input_checksum_ack;
  assign input_eth_rx_ack = s_input_eth_rx_ack;
  assign input_rs232_rx_ack = s_input_rs232_rx_ack;
  assign output_checksum_stb = s_output_checksum_stb;
  assign output_checksum = s_output_checksum;
  assign output_leds_stb = s_output_leds_stb;
  assign output_leds = s_output_leds;
  assign output_eth_tx_stb = s_output_eth_tx_stb;
  assign output_eth_tx = s_output_eth_tx;
  assign output_rs232_tx_stb = s_output_rs232_tx_stb;
  assign output_rs232_tx = s_output_rs232_tx;

endmodule
